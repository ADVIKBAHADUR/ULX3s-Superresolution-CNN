module modelReader(input wire clk,          // Clock
    input wire rst_n,        // Reset (active low)
    output reg [31:0] Weights [0:4][0:63][0:63][0:2][0:2], reg signed [31:0] Biases[0:4][0:63]);


// 5D Register to store convolution weights: [ConvLayer][Kernel][Depth][Height][Width]
// Fixed-point format: 16 fractional bits
reg signed [31:0] conv_weights[0:4][0:63][0:63][0:2][0:2] = '{
// Weights for conv1_weight
{
{
{{15'sd8400, 15'sd-12340, 13'sd3527}, {15'sd-12066, 15'sd-11606, 13'sd-2983}, {14'sd5793, 14'sd4791, 14'sd6601}},
{{14'sd-4491, 12'sd1269, 13'sd3175}, {14'sd4569, 15'sd-9277, 12'sd-1853}, {14'sd7041, 15'sd10070, 15'sd-10451}},
{{15'sd9065, 14'sd4972, 15'sd8974}, {13'sd-2049, 13'sd2351, 15'sd-9675}, {13'sd-2470, 15'sd13758, 13'sd3394}}},
{
{{14'sd6521, 14'sd6441, 12'sd1938}, {13'sd3792, 14'sd7267, 15'sd8900}, {12'sd1063, 13'sd-2078, 13'sd-3476}},
{{14'sd-6434, 14'sd-5689, 12'sd1211}, {15'sd11563, 15'sd12513, 14'sd-4893}, {15'sd13114, 15'sd10153, 13'sd-4040}},
{{15'sd-9517, 15'sd8371, 14'sd-4571}, {15'sd12415, 15'sd8479, 14'sd7376}, {14'sd5703, 15'sd-9070, 15'sd-11924}}},
{
{{15'sd11783, 15'sd-8289, 15'sd8968}, {14'sd5811, 15'sd-12238, 11'sd-922}, {14'sd7923, 14'sd-5686, 14'sd5332}},
{{13'sd3409, 13'sd-3990, 14'sd-8072}, {14'sd-4483, 14'sd-7349, 14'sd6119}, {14'sd-4164, 15'sd12792, 14'sd4533}},
{{15'sd-10004, 11'sd-579, 15'sd-11805}, {14'sd-7267, 13'sd2492, 13'sd3858}, {15'sd-10967, 15'sd8647, 15'sd-12127}}},
{
{{15'sd11858, 14'sd-6996, 14'sd7224}, {14'sd-7001, 14'sd-5333, 14'sd4204}, {13'sd-2151, 15'sd-8662, 12'sd2042}},
{{15'sd8727, 13'sd2976, 15'sd-13083}, {14'sd6794, 13'sd3909, 13'sd-2834}, {15'sd-11710, 14'sd-4380, 15'sd-11136}},
{{12'sd-2046, 14'sd-5336, 15'sd-9768}, {12'sd-1944, 15'sd-11460, 12'sd1240}, {15'sd-13891, 15'sd8944, 15'sd-9573}}},
{
{{14'sd-6883, 14'sd4154, 14'sd4515}, {11'sd522, 15'sd11772, 10'sd384}, {12'sd-1184, 13'sd4066, 12'sd1309}},
{{14'sd-6023, 15'sd-12426, 15'sd-9715}, {12'sd-1533, 13'sd-2148, 9'sd-197}, {14'sd-6352, 13'sd-2916, 14'sd-4353}},
{{13'sd-4035, 15'sd-11078, 13'sd3422}, {14'sd-4350, 14'sd5432, 14'sd-4991}, {15'sd9413, 13'sd3690, 15'sd10133}}},
{
{{15'sd-13284, 15'sd8662, 15'sd-10225}, {14'sd-7042, 14'sd-5808, 11'sd-978}, {15'sd9728, 14'sd-4305, 10'sd-504}},
{{14'sd-8125, 14'sd-6150, 12'sd-1318}, {13'sd2175, 15'sd9235, 12'sd-1260}, {15'sd11559, 14'sd4584, 15'sd-11739}},
{{15'sd14582, 15'sd11355, 15'sd-14167}, {14'sd-8059, 13'sd3812, 14'sd-6259}, {15'sd8639, 13'sd-2422, 15'sd-8737}}},
{
{{13'sd-4037, 15'sd10739, 8'sd120}, {15'sd-11372, 6'sd19, 14'sd-7235}, {13'sd3014, 10'sd-504, 13'sd2941}},
{{14'sd-5731, 14'sd7332, 13'sd3036}, {14'sd7995, 12'sd-1309, 15'sd-10295}, {14'sd-5714, 13'sd3004, 15'sd-13384}},
{{14'sd-5551, 13'sd-3157, 15'sd10471}, {15'sd10565, 15'sd-10152, 15'sd-9800}, {11'sd-652, 15'sd-13361, 13'sd-3955}}},
{
{{13'sd-2455, 15'sd-11059, 14'sd7836}, {14'sd6878, 15'sd8787, 14'sd-6433}, {10'sd500, 12'sd-1430, 13'sd-3214}},
{{13'sd2632, 14'sd5869, 15'sd-11575}, {14'sd7268, 15'sd9687, 11'sd895}, {10'sd436, 14'sd-4505, 15'sd-13128}},
{{15'sd9559, 15'sd-16043, 15'sd-14653}, {14'sd-4492, 7'sd-52, 15'sd-15591}, {14'sd4852, 13'sd-4041, 13'sd-2959}}},
{
{{15'sd9856, 15'sd11006, 14'sd4439}, {14'sd-7019, 14'sd-5085, 12'sd-1850}, {15'sd-10526, 14'sd5803, 15'sd11622}},
{{13'sd3478, 13'sd2287, 15'sd-8919}, {15'sd-11723, 14'sd-5744, 13'sd2651}, {14'sd5634, 13'sd3760, 15'sd12852}},
{{15'sd13781, 14'sd-7903, 15'sd13192}, {14'sd-4131, 10'sd348, 13'sd2151}, {15'sd8990, 9'sd164, 14'sd-7370}}},
{
{{15'sd11092, 15'sd-9618, 14'sd5862}, {15'sd9933, 13'sd2577, 14'sd-5507}, {12'sd1448, 12'sd1308, 15'sd9014}},
{{14'sd6012, 15'sd-13573, 14'sd5395}, {12'sd-1698, 15'sd8268, 13'sd-2552}, {15'sd-12822, 15'sd-12715, 14'sd-6609}},
{{15'sd10062, 15'sd-9977, 11'sd-753}, {15'sd10962, 13'sd3509, 15'sd-12891}, {14'sd-7801, 12'sd-1604, 14'sd-6488}}},
{
{{13'sd2524, 14'sd6314, 12'sd-1739}, {14'sd4872, 15'sd-11695, 14'sd-5754}, {15'sd8222, 15'sd-8660, 15'sd8372}},
{{12'sd1378, 15'sd-9370, 14'sd4397}, {13'sd3507, 14'sd6810, 14'sd4272}, {12'sd-1225, 11'sd-764, 14'sd-4117}},
{{14'sd-7172, 15'sd-14237, 14'sd-4231}, {13'sd-4043, 14'sd6554, 15'sd-11905}, {15'sd-13797, 14'sd-4559, 15'sd8778}}},
{
{{12'sd-1106, 15'sd-11811, 14'sd4909}, {12'sd1350, 14'sd-7235, 13'sd3618}, {12'sd1504, 8'sd126, 11'sd-965}},
{{15'sd-10316, 15'sd-11370, 15'sd-11020}, {12'sd-2040, 15'sd10409, 14'sd6328}, {13'sd2410, 15'sd11920, 14'sd7433}},
{{15'sd-10860, 15'sd8785, 14'sd6390}, {11'sd519, 13'sd3984, 13'sd-2844}, {15'sd12786, 15'sd9716, 15'sd10781}}},
{
{{13'sd4084, 15'sd12240, 15'sd10956}, {14'sd7864, 14'sd-6895, 15'sd10433}, {15'sd9043, 14'sd6826, 15'sd13181}},
{{15'sd11863, 12'sd2019, 13'sd3597}, {12'sd-1098, 14'sd5620, 15'sd-11482}, {15'sd-10095, 12'sd1504, 15'sd-11558}},
{{14'sd5875, 12'sd1407, 14'sd4321}, {15'sd-10813, 13'sd3150, 15'sd12744}, {14'sd-5093, 14'sd-6562, 15'sd-11046}}},
{
{{14'sd4175, 12'sd1835, 9'sd-153}, {14'sd5391, 13'sd-2082, 15'sd8381}, {13'sd-2965, 13'sd-2743, 14'sd-6579}},
{{15'sd9921, 15'sd-9833, 14'sd-6692}, {13'sd3987, 14'sd-5961, 14'sd4770}, {13'sd-3618, 12'sd-1427, 15'sd11977}},
{{14'sd-5243, 15'sd-13693, 15'sd-8793}, {15'sd-10975, 13'sd-2819, 13'sd3916}, {14'sd6189, 10'sd-495, 15'sd11892}}},
{
{{13'sd-2568, 14'sd-8104, 15'sd-11033}, {14'sd6213, 12'sd-1773, 14'sd7658}, {15'sd-12706, 14'sd-4829, 15'sd-11976}},
{{15'sd-8707, 14'sd4394, 15'sd-10868}, {11'sd-686, 15'sd-12256, 14'sd-5643}, {15'sd-14423, 15'sd-9606, 12'sd-1740}},
{{15'sd-14131, 13'sd-3607, 15'sd9424}, {11'sd870, 14'sd-7143, 15'sd9416}, {14'sd-4179, 15'sd9795, 14'sd5942}}},
{
{{11'sd-513, 15'sd12201, 15'sd10235}, {15'sd9958, 14'sd-6661, 15'sd10851}, {14'sd5779, 15'sd10431, 10'sd494}},
{{14'sd6396, 15'sd-9045, 13'sd-3160}, {14'sd5659, 15'sd12405, 13'sd-2167}, {14'sd-4370, 15'sd12471, 14'sd4365}},
{{14'sd7389, 15'sd9504, 15'sd11083}, {15'sd-12227, 12'sd-1808, 4'sd4}, {14'sd-4142, 15'sd-9812, 15'sd11957}}},
{
{{15'sd10251, 15'sd-9846, 14'sd-6483}, {13'sd3109, 13'sd-2295, 13'sd-4092}, {11'sd-514, 12'sd-1287, 12'sd1050}},
{{14'sd4352, 15'sd-10238, 12'sd1290}, {13'sd2967, 15'sd9457, 14'sd-5014}, {13'sd3956, 15'sd8220, 14'sd4689}},
{{11'sd771, 15'sd11178, 13'sd2771}, {15'sd-11516, 15'sd10430, 14'sd-7564}, {15'sd11936, 14'sd7056, 11'sd-662}}},
{
{{15'sd10292, 9'sd-211, 13'sd2375}, {14'sd-6564, 15'sd13262, 15'sd9192}, {12'sd-1178, 13'sd-2055, 14'sd5155}},
{{15'sd-9184, 15'sd-13037, 6'sd17}, {12'sd1136, 12'sd-1924, 15'sd-13006}, {15'sd-12654, 14'sd4629, 11'sd-595}},
{{14'sd-6667, 14'sd5495, 14'sd-7148}, {12'sd1079, 14'sd-7284, 14'sd6845}, {15'sd-13418, 14'sd7325, 14'sd-7005}}},
{
{{14'sd5126, 14'sd-6791, 12'sd1525}, {15'sd8789, 14'sd4201, 13'sd2651}, {14'sd-7997, 15'sd-9856, 15'sd-10930}},
{{14'sd-7269, 7'sd-42, 14'sd7544}, {15'sd9526, 14'sd4699, 13'sd-4021}, {15'sd-13175, 13'sd-2406, 14'sd-5790}},
{{12'sd1306, 14'sd7538, 14'sd-6723}, {15'sd-10206, 12'sd-1235, 15'sd9735}, {12'sd-1086, 14'sd-5582, 15'sd-10234}}},
{
{{13'sd3028, 11'sd725, 13'sd-2203}, {15'sd-8585, 15'sd-8787, 15'sd-9311}, {15'sd-10522, 14'sd-5578, 14'sd-5461}},
{{15'sd11823, 15'sd-9888, 14'sd6888}, {14'sd-4578, 14'sd5988, 15'sd-11578}, {13'sd3010, 15'sd9198, 14'sd4384}},
{{15'sd12840, 15'sd8333, 14'sd-6200}, {14'sd-7800, 11'sd740, 15'sd8452}, {15'sd11117, 14'sd-6993, 14'sd5244}}},
{
{{15'sd-12710, 13'sd-2729, 15'sd-10561}, {15'sd-12480, 15'sd11590, 15'sd-9810}, {14'sd6433, 14'sd-4108, 14'sd4191}},
{{14'sd-6865, 14'sd6416, 14'sd7453}, {14'sd6498, 12'sd-1650, 15'sd-12608}, {14'sd-4507, 13'sd-2295, 14'sd-7184}},
{{14'sd-6990, 11'sd877, 14'sd-4488}, {14'sd-6427, 14'sd7825, 11'sd564}, {7'sd-46, 13'sd3794, 12'sd1873}}},
{
{{13'sd-3363, 14'sd-5555, 14'sd7166}, {14'sd7860, 11'sd-892, 14'sd-7355}, {12'sd1414, 14'sd7781, 11'sd847}},
{{15'sd8625, 14'sd6866, 12'sd-1355}, {14'sd-5383, 14'sd7780, 14'sd5693}, {15'sd9902, 13'sd-3830, 15'sd-10876}},
{{13'sd3266, 15'sd12835, 13'sd-3716}, {14'sd-5977, 14'sd7845, 14'sd5210}, {15'sd13652, 15'sd11808, 13'sd2244}}},
{
{{15'sd9076, 15'sd-10498, 14'sd-8008}, {15'sd10881, 15'sd13698, 14'sd5564}, {14'sd7474, 15'sd8289, 15'sd11155}},
{{14'sd-6946, 11'sd589, 14'sd-7765}, {13'sd-3626, 14'sd7923, 13'sd4078}, {12'sd-1161, 13'sd2791, 13'sd-4094}},
{{15'sd8391, 14'sd-5526, 15'sd10640}, {15'sd-9060, 15'sd9522, 15'sd8434}, {15'sd10893, 13'sd2292, 13'sd-3964}}},
{
{{8'sd-76, 14'sd6869, 15'sd-10054}, {14'sd-5153, 15'sd10750, 12'sd-1962}, {14'sd-6766, 13'sd-2054, 13'sd3985}},
{{13'sd3367, 15'sd8380, 11'sd786}, {13'sd-3298, 13'sd3947, 15'sd11398}, {15'sd-12603, 15'sd-10261, 15'sd10069}},
{{13'sd2356, 14'sd5241, 14'sd4710}, {14'sd7491, 14'sd-4406, 13'sd2730}, {15'sd-10913, 15'sd-9898, 11'sd-936}}},
{
{{14'sd5514, 11'sd518, 15'sd-9585}, {6'sd27, 15'sd9250, 14'sd5493}, {15'sd11158, 13'sd3459, 14'sd-7738}},
{{13'sd2595, 14'sd5405, 14'sd4581}, {15'sd-8874, 13'sd-3277, 14'sd-7495}, {15'sd9496, 14'sd4656, 13'sd-3865}},
{{13'sd3186, 14'sd7223, 11'sd564}, {15'sd-10385, 14'sd-6503, 15'sd-9051}, {14'sd-6164, 12'sd-1405, 12'sd-1537}}},
{
{{14'sd-4360, 13'sd-2572, 13'sd2321}, {15'sd10529, 13'sd4034, 13'sd2487}, {15'sd10532, 14'sd6241, 15'sd12567}},
{{15'sd-12109, 12'sd-1493, 15'sd-9675}, {12'sd1084, 13'sd-2188, 15'sd-12490}, {14'sd-5427, 14'sd5185, 14'sd6016}},
{{15'sd-12303, 14'sd6373, 14'sd-4858}, {15'sd-12419, 9'sd160, 12'sd1504}, {14'sd-6123, 14'sd4233, 15'sd-11872}}},
{
{{13'sd-2610, 15'sd13760, 15'sd-10165}, {12'sd1613, 12'sd-2000, 15'sd8940}, {15'sd-12456, 15'sd11545, 14'sd5035}},
{{15'sd10679, 14'sd-5011, 15'sd8553}, {15'sd8994, 11'sd-946, 13'sd-2735}, {10'sd-413, 14'sd7922, 15'sd12052}},
{{15'sd-12458, 14'sd-5796, 15'sd-13172}, {16'sd-17613, 15'sd-11078, 14'sd-7023}, {16'sd-19290, 14'sd-6731, 10'sd476}}},
{
{{14'sd-5153, 15'sd-11653, 9'sd168}, {15'sd-10734, 14'sd-7370, 13'sd-2173}, {13'sd-2358, 13'sd-4014, 12'sd1676}},
{{14'sd-6894, 15'sd-10705, 14'sd-5346}, {15'sd-9284, 14'sd-5633, 14'sd-5599}, {15'sd-11593, 14'sd-4790, 15'sd-11739}},
{{12'sd-1711, 15'sd8965, 14'sd7217}, {14'sd-8184, 15'sd-12772, 15'sd8742}, {12'sd1402, 11'sd1000, 15'sd9959}}},
{
{{14'sd6515, 14'sd-4384, 15'sd-11305}, {13'sd2546, 13'sd-2183, 15'sd-13325}, {14'sd5884, 14'sd5953, 14'sd-6022}},
{{14'sd-6677, 12'sd-1307, 12'sd1624}, {13'sd3823, 13'sd2571, 13'sd4059}, {13'sd-2178, 15'sd-8471, 13'sd-3783}},
{{15'sd-13238, 14'sd-5883, 13'sd2359}, {15'sd-9078, 12'sd1800, 13'sd3350}, {14'sd-5703, 11'sd-818, 14'sd7080}}},
{
{{13'sd-4055, 14'sd7665, 15'sd9601}, {15'sd-12173, 13'sd-2528, 13'sd-3700}, {14'sd-7215, 12'sd-1102, 12'sd1884}},
{{12'sd1144, 11'sd686, 15'sd14302}, {14'sd-6833, 15'sd10292, 15'sd12731}, {14'sd7341, 14'sd-6452, 15'sd8197}},
{{14'sd7150, 13'sd-2735, 13'sd-3877}, {15'sd-12717, 15'sd-12358, 12'sd1978}, {14'sd-6931, 7'sd-49, 14'sd-4482}}},
{
{{14'sd-7430, 14'sd5355, 15'sd-10026}, {13'sd-3321, 15'sd10681, 13'sd3813}, {13'sd2493, 13'sd3671, 12'sd1777}},
{{13'sd-3937, 14'sd7251, 12'sd1152}, {12'sd-1615, 13'sd2820, 14'sd6146}, {13'sd3746, 15'sd-9531, 12'sd1754}},
{{15'sd-9829, 15'sd11698, 15'sd-8822}, {13'sd2529, 15'sd11699, 13'sd-2620}, {15'sd13836, 15'sd10387, 15'sd-9649}}},
{
{{12'sd-1977, 11'sd528, 15'sd-9164}, {15'sd10663, 12'sd1024, 15'sd-11349}, {12'sd-1724, 13'sd2865, 14'sd4376}},
{{10'sd326, 15'sd12050, 15'sd-10461}, {12'sd1997, 14'sd4423, 13'sd2881}, {14'sd6940, 15'sd-9212, 14'sd4460}},
{{15'sd-11049, 12'sd-1373, 15'sd12620}, {15'sd10527, 13'sd4044, 14'sd5746}, {10'sd469, 15'sd-11705, 15'sd10365}}},
{
{{15'sd-11559, 15'sd9928, 15'sd11229}, {14'sd-7860, 15'sd-9572, 15'sd-9303}, {12'sd-1925, 15'sd9064, 15'sd11561}},
{{14'sd4786, 15'sd-12675, 14'sd6698}, {14'sd4250, 14'sd5074, 14'sd5011}, {13'sd-2748, 12'sd-1865, 12'sd-1567}},
{{15'sd-9175, 15'sd10886, 15'sd11872}, {10'sd426, 15'sd9581, 12'sd-1083}, {13'sd-3336, 14'sd6931, 15'sd11246}}},
{
{{13'sd3877, 14'sd7228, 15'sd10435}, {12'sd-1446, 15'sd-8713, 15'sd-11942}, {14'sd-6643, 15'sd-11099, 15'sd-12483}},
{{15'sd-11726, 15'sd12337, 14'sd-4119}, {15'sd-9670, 15'sd-9830, 15'sd12053}, {12'sd1164, 12'sd1359, 14'sd4355}},
{{13'sd3219, 13'sd-4078, 15'sd14123}, {13'sd2488, 12'sd1088, 15'sd10983}, {14'sd4464, 12'sd1361, 13'sd3824}}},
{
{{15'sd-10413, 13'sd2688, 13'sd2865}, {14'sd-4575, 15'sd-12102, 15'sd10529}, {14'sd6452, 15'sd-10452, 14'sd4556}},
{{15'sd-13089, 15'sd-9080, 15'sd10424}, {15'sd9656, 15'sd8910, 11'sd-931}, {13'sd2725, 15'sd8294, 12'sd1118}},
{{14'sd-6220, 15'sd-8903, 15'sd9675}, {13'sd3458, 15'sd11303, 13'sd-2158}, {13'sd2086, 14'sd4118, 15'sd8397}}},
{
{{14'sd7380, 15'sd-11720, 15'sd-9287}, {14'sd-7765, 12'sd-1775, 13'sd2983}, {14'sd7434, 14'sd-4470, 12'sd1723}},
{{14'sd4271, 14'sd-7525, 15'sd-12206}, {13'sd2548, 15'sd11163, 14'sd4943}, {11'sd529, 15'sd-9181, 14'sd-4664}},
{{14'sd7757, 15'sd9927, 13'sd-2642}, {12'sd-1685, 14'sd-6596, 14'sd-6940}, {15'sd-10664, 14'sd-5809, 13'sd2276}}},
{
{{15'sd-8589, 13'sd-2654, 13'sd-3768}, {14'sd-6240, 13'sd-2997, 15'sd-9932}, {14'sd-6542, 13'sd-2239, 14'sd5247}},
{{14'sd4366, 15'sd12105, 11'sd636}, {15'sd10313, 14'sd-4300, 12'sd-1394}, {15'sd8329, 15'sd10109, 13'sd-3081}},
{{12'sd1720, 15'sd8708, 12'sd-1545}, {14'sd-5936, 14'sd-6510, 12'sd1980}, {13'sd-3570, 14'sd-7314, 15'sd12712}}},
{
{{14'sd-5338, 14'sd7580, 13'sd3954}, {14'sd-6902, 14'sd-4328, 14'sd7805}, {14'sd5701, 14'sd4752, 13'sd2594}},
{{14'sd-5182, 14'sd-5645, 9'sd-193}, {13'sd3268, 15'sd-11348, 14'sd-7876}, {13'sd-2590, 13'sd3903, 11'sd-722}},
{{15'sd8796, 15'sd-11858, 13'sd2353}, {14'sd6241, 14'sd-6538, 15'sd-10607}, {15'sd-10344, 14'sd-6698, 12'sd1803}}},
{
{{13'sd-3654, 14'sd-6198, 15'sd-11061}, {14'sd-6242, 12'sd-1078, 15'sd8559}, {14'sd4675, 9'sd175, 15'sd10746}},
{{15'sd-12142, 15'sd-8220, 14'sd8117}, {15'sd9832, 13'sd4072, 11'sd-658}, {10'sd-463, 7'sd50, 13'sd-2338}},
{{12'sd-1934, 15'sd-10441, 15'sd-15527}, {15'sd-11475, 15'sd8267, 11'sd-772}, {13'sd-4094, 13'sd-3304, 13'sd-3604}}},
{
{{15'sd10736, 15'sd-10956, 14'sd6842}, {13'sd-2117, 15'sd-9821, 15'sd12275}, {12'sd1763, 14'sd7787, 13'sd3982}},
{{14'sd6076, 12'sd1668, 15'sd-10835}, {15'sd-11194, 14'sd-7935, 14'sd-4496}, {14'sd4447, 13'sd-3370, 15'sd8726}},
{{14'sd7045, 15'sd8650, 13'sd-3736}, {15'sd13592, 15'sd-8947, 15'sd10119}, {13'sd-2892, 10'sd-413, 14'sd-7404}}},
{
{{12'sd-1308, 13'sd-2513, 14'sd7950}, {14'sd-7456, 13'sd3605, 15'sd9038}, {15'sd-9386, 13'sd3376, 14'sd5189}},
{{15'sd-8373, 15'sd-10741, 13'sd-3724}, {15'sd10184, 14'sd-6300, 12'sd1937}, {15'sd9238, 15'sd-13045, 15'sd-11467}},
{{15'sd10751, 15'sd-9762, 15'sd9605}, {15'sd8491, 7'sd44, 15'sd-12601}, {11'sd-841, 15'sd-8434, 15'sd-11760}}},
{
{{15'sd-11085, 15'sd-11148, 15'sd10160}, {15'sd8199, 13'sd-2128, 14'sd-5338}, {15'sd11293, 15'sd11863, 15'sd11297}},
{{14'sd-4800, 15'sd-10610, 14'sd8027}, {13'sd-2088, 14'sd4330, 14'sd-4874}, {12'sd-1785, 14'sd-5488, 14'sd5035}},
{{14'sd-6046, 14'sd-6610, 9'sd245}, {15'sd11117, 11'sd-790, 14'sd7956}, {14'sd-7760, 12'sd1042, 14'sd-4284}}},
{
{{15'sd-9950, 14'sd-5018, 9'sd145}, {15'sd10100, 14'sd-6284, 13'sd-3687}, {14'sd5935, 15'sd-10779, 14'sd4999}},
{{15'sd-8888, 14'sd6951, 15'sd9301}, {13'sd-4044, 12'sd1304, 13'sd3984}, {15'sd-9094, 11'sd-538, 15'sd-9055}},
{{14'sd-6786, 15'sd-10925, 14'sd-8093}, {15'sd-15428, 15'sd-14735, 15'sd9145}, {15'sd-8868, 13'sd2700, 14'sd-4494}}},
{
{{14'sd-7239, 14'sd-5810, 14'sd6161}, {13'sd3142, 14'sd6479, 10'sd-403}, {15'sd15077, 14'sd5427, 10'sd431}},
{{12'sd1363, 12'sd-1286, 14'sd-6093}, {13'sd3905, 15'sd8978, 15'sd-9748}, {15'sd10201, 10'sd379, 14'sd7019}},
{{15'sd-11031, 15'sd-14852, 15'sd-9962}, {15'sd-12660, 15'sd9904, 14'sd-5268}, {12'sd1614, 14'sd-5517, 15'sd10604}}},
{
{{14'sd5500, 12'sd-1736, 15'sd9767}, {13'sd-3756, 14'sd5183, 14'sd-6369}, {15'sd-10731, 13'sd3895, 10'sd487}},
{{13'sd2882, 14'sd8191, 14'sd-5555}, {11'sd-781, 15'sd10552, 15'sd-10475}, {9'sd188, 14'sd7114, 12'sd-1439}},
{{12'sd1222, 14'sd7363, 15'sd10110}, {12'sd1151, 15'sd-10021, 12'sd-1525}, {15'sd-13739, 12'sd-1388, 9'sd233}}},
{
{{15'sd-8430, 15'sd-10005, 11'sd946}, {7'sd-58, 15'sd9576, 14'sd-4833}, {13'sd2374, 11'sd-968, 15'sd8647}},
{{15'sd-10929, 15'sd12264, 15'sd-12397}, {15'sd11641, 15'sd10473, 15'sd-9348}, {13'sd-2390, 14'sd7999, 15'sd8716}},
{{8'sd82, 14'sd6073, 14'sd-6149}, {7'sd-51, 14'sd7885, 12'sd1408}, {15'sd13692, 12'sd1296, 13'sd-3404}}},
{
{{13'sd2238, 13'sd-3011, 10'sd510}, {14'sd-6196, 14'sd7043, 12'sd-1407}, {15'sd-12674, 8'sd-78, 14'sd5477}},
{{13'sd-2852, 14'sd7696, 10'sd404}, {15'sd12581, 15'sd10710, 14'sd5707}, {12'sd1249, 14'sd8092, 14'sd-6006}},
{{13'sd-3611, 14'sd4256, 14'sd7387}, {14'sd-8008, 15'sd11848, 15'sd11624}, {15'sd-12169, 15'sd-10205, 14'sd4643}}},
{
{{3'sd3, 14'sd-7182, 15'sd11746}, {15'sd-9656, 14'sd7647, 11'sd1023}, {15'sd-11311, 13'sd2317, 14'sd8018}},
{{13'sd-2340, 15'sd-8426, 12'sd-1852}, {13'sd3612, 14'sd-6231, 13'sd-3945}, {14'sd-8093, 14'sd-4549, 15'sd11968}},
{{14'sd-7927, 15'sd-10945, 15'sd11427}, {15'sd-14683, 15'sd-8999, 12'sd-1318}, {14'sd5015, 14'sd-5285, 14'sd5660}}},
{
{{15'sd-9319, 14'sd-7244, 13'sd-3743}, {15'sd-11118, 14'sd6090, 15'sd-13717}, {15'sd-10018, 15'sd-14183, 15'sd-11393}},
{{15'sd-8212, 15'sd8621, 14'sd-6786}, {14'sd6933, 12'sd1495, 14'sd8143}, {14'sd-7519, 15'sd13041, 12'sd-1381}},
{{13'sd2857, 15'sd-11902, 15'sd-14057}, {13'sd-2925, 15'sd10008, 15'sd-13108}, {14'sd-5742, 14'sd-7839, 15'sd-13687}}},
{
{{10'sd500, 15'sd10958, 15'sd-11958}, {15'sd-9601, 14'sd7536, 15'sd10695}, {14'sd-5180, 13'sd4073, 14'sd-7167}},
{{11'sd590, 14'sd7956, 15'sd9650}, {12'sd-1445, 12'sd1091, 14'sd-5382}, {13'sd-2515, 12'sd-1105, 14'sd7510}},
{{13'sd3606, 15'sd9216, 14'sd6206}, {12'sd-1367, 15'sd13318, 15'sd8350}, {13'sd3196, 15'sd14205, 14'sd-4292}}},
{
{{13'sd3761, 15'sd9462, 13'sd-3472}, {14'sd-5325, 13'sd-2533, 14'sd5662}, {12'sd-1140, 11'sd-784, 12'sd1208}},
{{15'sd-14421, 15'sd-13942, 14'sd5998}, {14'sd6454, 14'sd-6274, 14'sd4823}, {13'sd-3352, 15'sd-12713, 15'sd9748}},
{{14'sd-6713, 12'sd1457, 15'sd13400}, {14'sd8122, 14'sd-5328, 13'sd-3471}, {12'sd-1047, 12'sd1783, 15'sd11062}}},
{
{{14'sd7103, 12'sd1247, 9'sd-191}, {13'sd-3332, 15'sd-12051, 13'sd-2330}, {14'sd5189, 15'sd12326, 15'sd-9780}},
{{14'sd5150, 14'sd-4141, 14'sd6877}, {13'sd-2725, 15'sd11830, 14'sd5338}, {14'sd-7722, 15'sd9449, 15'sd-10265}},
{{14'sd4132, 14'sd-7448, 14'sd-7898}, {10'sd272, 15'sd10982, 14'sd-5226}, {15'sd14282, 13'sd2425, 13'sd-2458}}},
{
{{15'sd-10382, 15'sd-9965, 13'sd2452}, {15'sd11027, 15'sd-9215, 14'sd-4130}, {15'sd8200, 14'sd-4123, 14'sd-4580}},
{{11'sd-593, 13'sd-2764, 13'sd3450}, {13'sd3047, 15'sd-8877, 13'sd2813}, {15'sd-12656, 14'sd-4541, 14'sd-7546}},
{{14'sd-4319, 14'sd5913, 8'sd-126}, {13'sd2331, 14'sd-4810, 14'sd-4352}, {15'sd9985, 8'sd-81, 14'sd8174}}},
{
{{13'sd-2059, 13'sd-3602, 11'sd-934}, {15'sd9029, 15'sd-9152, 15'sd13005}, {15'sd8264, 13'sd3021, 13'sd3214}},
{{10'sd325, 15'sd9884, 10'sd340}, {14'sd-6097, 14'sd5477, 15'sd-9636}, {8'sd70, 14'sd5368, 14'sd7913}},
{{15'sd8378, 14'sd-5872, 15'sd-10771}, {15'sd-10686, 15'sd-13027, 15'sd11889}, {15'sd-12091, 15'sd-13009, 13'sd-2951}}},
{
{{13'sd-3824, 13'sd3956, 14'sd-5079}, {14'sd-5636, 14'sd5848, 15'sd12073}, {12'sd-1697, 12'sd1451, 15'sd12628}},
{{13'sd2319, 14'sd-4336, 13'sd3582}, {13'sd2180, 14'sd-4725, 12'sd-2035}, {15'sd-12368, 14'sd-5120, 13'sd-3810}},
{{14'sd-7059, 15'sd9490, 14'sd5021}, {13'sd-2550, 11'sd887, 15'sd-11326}, {15'sd-10752, 15'sd-11901, 13'sd-4052}}},
{
{{15'sd-9651, 15'sd-8851, 15'sd-10283}, {14'sd-6857, 14'sd-7807, 12'sd2030}, {14'sd-4666, 14'sd7627, 13'sd-2900}},
{{15'sd9390, 15'sd9158, 14'sd6188}, {11'sd-884, 15'sd11282, 13'sd-3753}, {14'sd4935, 12'sd-1261, 14'sd-7309}},
{{15'sd9770, 15'sd9026, 14'sd5412}, {13'sd3283, 15'sd-11582, 15'sd-12008}, {13'sd3532, 15'sd11498, 9'sd-181}}},
{
{{14'sd6110, 13'sd3290, 14'sd4394}, {14'sd-4432, 13'sd-2066, 15'sd8756}, {12'sd-1688, 15'sd9734, 14'sd5074}},
{{15'sd11360, 14'sd-6323, 14'sd5802}, {12'sd-1131, 15'sd-9193, 10'sd-429}, {15'sd-11594, 14'sd-6656, 8'sd115}},
{{13'sd-2787, 15'sd-10626, 14'sd7444}, {11'sd902, 14'sd-6348, 12'sd-1290}, {15'sd11827, 6'sd-16, 15'sd8755}}},
{
{{13'sd3469, 12'sd1927, 15'sd12807}, {14'sd-4849, 13'sd4009, 15'sd11249}, {13'sd3503, 15'sd-10057, 14'sd-4488}},
{{14'sd-7690, 14'sd-7483, 15'sd-9902}, {15'sd11423, 14'sd4704, 14'sd-7305}, {14'sd-5552, 14'sd-6505, 15'sd9134}},
{{14'sd7106, 14'sd-7865, 13'sd4021}, {11'sd-1021, 14'sd5592, 15'sd12072}, {13'sd2500, 14'sd4941, 15'sd-12617}}},
{
{{6'sd-25, 13'sd-2847, 10'sd-371}, {13'sd-3079, 15'sd-10544, 13'sd3709}, {15'sd10987, 11'sd844, 15'sd11231}},
{{15'sd-11288, 15'sd-8938, 15'sd-10762}, {14'sd-7471, 13'sd2790, 15'sd-8846}, {14'sd-5585, 14'sd4644, 14'sd-7623}},
{{13'sd3089, 13'sd-3443, 14'sd-5407}, {13'sd-2054, 15'sd-12783, 14'sd-7530}, {13'sd-2779, 13'sd-2829, 15'sd-12405}}},
{
{{15'sd9983, 12'sd1514, 15'sd-9114}, {15'sd-12427, 15'sd-11696, 11'sd-769}, {15'sd-14941, 15'sd11645, 14'sd5656}},
{{15'sd-12229, 13'sd-3181, 14'sd-4128}, {14'sd-6781, 11'sd961, 13'sd3855}, {13'sd2577, 15'sd10338, 13'sd-2985}},
{{13'sd2351, 14'sd7119, 15'sd9617}, {15'sd-10193, 11'sd-817, 15'sd10425}, {15'sd-13954, 15'sd-9070, 15'sd-12239}}},
{
{{13'sd-3819, 14'sd6642, 15'sd10949}, {15'sd-10021, 15'sd8987, 15'sd9761}, {14'sd-5621, 13'sd3426, 15'sd-10817}},
{{14'sd6706, 15'sd-9378, 15'sd-12956}, {13'sd-2708, 15'sd-11197, 15'sd8842}, {14'sd-4959, 14'sd6339, 12'sd-1323}},
{{14'sd5107, 15'sd13435, 11'sd-819}, {15'sd8909, 11'sd-958, 15'sd9569}, {14'sd7536, 14'sd6266, 15'sd13725}}},
{
{{13'sd2073, 14'sd-6831, 12'sd1420}, {14'sd6222, 13'sd3199, 14'sd-4720}, {13'sd-3537, 14'sd4806, 15'sd9949}},
{{14'sd-5155, 13'sd-3119, 13'sd-4063}, {14'sd7552, 15'sd9279, 14'sd5005}, {15'sd-10977, 15'sd-9110, 15'sd-12328}},
{{15'sd11607, 11'sd-735, 15'sd10118}, {13'sd-3455, 15'sd12099, 14'sd6370}, {15'sd-9137, 15'sd11643, 7'sd42}}},
{
{{14'sd-6955, 13'sd3107, 9'sd-229}, {14'sd-6183, 12'sd1732, 13'sd3687}, {15'sd-9189, 12'sd1143, 15'sd11434}},
{{15'sd10930, 15'sd-13228, 13'sd3526}, {15'sd11155, 14'sd5421, 15'sd-9279}, {14'sd5678, 11'sd-903, 10'sd-353}},
{{13'sd2802, 15'sd-9353, 15'sd-10188}, {14'sd-7417, 14'sd4714, 15'sd8797}, {11'sd919, 15'sd14446, 10'sd417}}},
{
{{13'sd-2132, 15'sd-12100, 15'sd-11288}, {15'sd12446, 14'sd-6618, 15'sd-13071}, {14'sd4903, 14'sd-7546, 15'sd-12967}},
{{15'sd10928, 13'sd3182, 15'sd-8717}, {15'sd-10306, 13'sd2501, 15'sd11528}, {14'sd-6154, 13'sd3670, 12'sd-1370}},
{{14'sd-5570, 14'sd-5980, 13'sd-3118}, {15'sd11119, 14'sd-6563, 15'sd-12524}, {14'sd-8129, 15'sd9292, 14'sd-7342}}}},
// Weights for conv2_weight
{
{
{{12'sd1250, 13'sd-2075, 13'sd2721}, {12'sd-1083, 12'sd1186, 11'sd-612}, {11'sd-846, 13'sd2334, 12'sd-1767}},
{{13'sd-2582, 12'sd1608, 13'sd2588}, {12'sd1671, 13'sd2446, 11'sd594}, {12'sd-1236, 11'sd876, 11'sd708}},
{{12'sd-1402, 12'sd-1586, 12'sd-1779}, {12'sd1789, 12'sd1227, 10'sd463}, {13'sd-2786, 8'sd77, 13'sd2300}},
{{12'sd1308, 13'sd-2148, 13'sd2481}, {11'sd877, 12'sd1999, 10'sd457}, {9'sd236, 11'sd791, 10'sd-360}},
{{13'sd3344, 12'sd1297, 11'sd619}, {12'sd1465, 13'sd2926, 14'sd4398}, {13'sd3355, 9'sd155, 13'sd3096}},
{{13'sd-2248, 12'sd1857, 10'sd339}, {13'sd-2326, 11'sd743, 13'sd-2587}, {12'sd1335, 10'sd415, 12'sd-1964}},
{{13'sd2550, 13'sd2155, 13'sd2654}, {13'sd3182, 13'sd-2159, 8'sd-117}, {12'sd1223, 11'sd817, 8'sd70}},
{{12'sd-1127, 13'sd2406, 10'sd-373}, {13'sd-2638, 11'sd-929, 13'sd2499}, {13'sd-2783, 11'sd-870, 10'sd-454}},
{{7'sd-61, 12'sd1348, 11'sd-759}, {11'sd875, 12'sd-1077, 10'sd460}, {12'sd2019, 13'sd-2154, 11'sd961}},
{{12'sd-1867, 13'sd2720, 12'sd1780}, {12'sd-1559, 11'sd893, 12'sd-1694}, {9'sd152, 9'sd128, 11'sd-704}},
{{11'sd-742, 13'sd-2428, 9'sd137}, {12'sd-1137, 11'sd659, 12'sd-1098}, {8'sd119, 11'sd975, 12'sd-1633}},
{{9'sd177, 13'sd-2884, 12'sd1197}, {13'sd-2072, 12'sd-1712, 10'sd296}, {13'sd2147, 13'sd2348, 11'sd593}},
{{13'sd2426, 8'sd78, 11'sd-1009}, {13'sd2743, 13'sd2991, 14'sd4494}, {11'sd-865, 11'sd550, 10'sd436}},
{{13'sd2065, 12'sd-1751, 12'sd1109}, {10'sd478, 13'sd-3153, 9'sd-178}, {12'sd-1197, 12'sd-1934, 12'sd-1995}},
{{12'sd-1989, 12'sd-1504, 13'sd-2913}, {13'sd-3380, 13'sd-2950, 12'sd1220}, {12'sd-1936, 8'sd-101, 13'sd2851}},
{{11'sd-570, 10'sd485, 12'sd1200}, {12'sd-1314, 12'sd-1472, 11'sd-809}, {9'sd224, 13'sd3150, 12'sd-1880}},
{{6'sd-28, 13'sd-2076, 12'sd1481}, {12'sd-1508, 11'sd-677, 12'sd1615}, {9'sd-224, 11'sd902, 12'sd1100}},
{{11'sd-595, 13'sd2113, 12'sd-1225}, {13'sd2419, 11'sd635, 9'sd-154}, {7'sd-59, 13'sd2632, 12'sd1617}},
{{11'sd934, 13'sd-2748, 11'sd959}, {12'sd-1499, 11'sd-596, 13'sd-3206}, {12'sd-1646, 12'sd-1345, 11'sd-980}},
{{13'sd2487, 13'sd-2094, 11'sd591}, {11'sd887, 12'sd-1665, 11'sd-568}, {10'sd-321, 13'sd-2736, 13'sd-3001}},
{{13'sd3079, 12'sd-1883, 11'sd-643}, {12'sd-1598, 11'sd932, 12'sd-1171}, {13'sd-2498, 11'sd-799, 11'sd-593}},
{{10'sd-426, 11'sd-931, 10'sd-454}, {9'sd162, 12'sd1336, 12'sd1133}, {9'sd227, 9'sd-146, 11'sd992}},
{{12'sd1138, 11'sd-676, 12'sd-1853}, {12'sd1298, 12'sd-1318, 6'sd29}, {10'sd413, 11'sd-656, 13'sd-2060}},
{{12'sd-1867, 13'sd2538, 13'sd2368}, {13'sd2341, 12'sd1415, 13'sd2259}, {13'sd-2232, 13'sd-2465, 11'sd651}},
{{12'sd1648, 12'sd1390, 12'sd1199}, {13'sd2490, 10'sd-342, 11'sd902}, {13'sd-2696, 12'sd-1831, 12'sd1352}},
{{13'sd-2248, 13'sd2110, 13'sd-2334}, {12'sd1744, 9'sd253, 12'sd1459}, {12'sd1512, 12'sd1525, 13'sd2384}},
{{12'sd-1693, 13'sd-2068, 12'sd-1910}, {12'sd1151, 13'sd-2480, 8'sd-106}, {12'sd-1049, 13'sd-4032, 11'sd1010}},
{{12'sd-1467, 12'sd1780, 12'sd-1451}, {12'sd-1800, 13'sd-2330, 12'sd1857}, {12'sd1594, 12'sd-1955, 13'sd-2243}},
{{13'sd-2907, 13'sd-3287, 10'sd346}, {13'sd-2123, 9'sd-129, 12'sd-1813}, {12'sd-1737, 13'sd-2339, 13'sd-2836}},
{{10'sd296, 13'sd-2117, 10'sd-446}, {10'sd428, 10'sd-403, 10'sd-436}, {9'sd136, 8'sd-103, 13'sd-2528}},
{{12'sd-1482, 12'sd1557, 11'sd-670}, {11'sd-815, 13'sd-2116, 11'sd794}, {12'sd1302, 11'sd-547, 10'sd490}},
{{12'sd1922, 13'sd-2548, 11'sd889}, {12'sd-1882, 12'sd-1160, 13'sd2445}, {13'sd-2063, 12'sd1986, 11'sd692}},
{{12'sd1265, 13'sd-2189, 10'sd495}, {12'sd1829, 10'sd-425, 12'sd-1105}, {13'sd2367, 11'sd-878, 13'sd-2535}},
{{8'sd73, 11'sd759, 12'sd1770}, {11'sd-747, 11'sd761, 12'sd-1430}, {12'sd-1567, 12'sd1040, 8'sd79}},
{{10'sd-445, 12'sd1680, 13'sd-3352}, {13'sd-2267, 12'sd-2005, 12'sd1134}, {13'sd2604, 13'sd-2206, 8'sd92}},
{{13'sd2351, 13'sd-2362, 12'sd1729}, {13'sd-2747, 12'sd-1194, 12'sd1311}, {12'sd1639, 13'sd-2499, 11'sd-896}},
{{13'sd2196, 12'sd-1370, 12'sd-1949}, {11'sd943, 13'sd-3730, 11'sd-744}, {12'sd-1162, 12'sd-1346, 14'sd-5518}},
{{11'sd808, 12'sd1894, 13'sd2251}, {12'sd1838, 12'sd-1526, 6'sd-22}, {11'sd-879, 10'sd359, 12'sd1922}},
{{11'sd-822, 12'sd1061, 9'sd177}, {12'sd-1918, 12'sd-1871, 12'sd-1209}, {12'sd1682, 12'sd1819, 12'sd-1848}},
{{12'sd-1506, 11'sd820, 12'sd-1564}, {13'sd2463, 9'sd222, 12'sd-1866}, {13'sd2758, 13'sd2084, 11'sd-1003}},
{{12'sd-1718, 13'sd2262, 14'sd4114}, {12'sd-1612, 11'sd719, 12'sd1604}, {12'sd-2029, 13'sd2911, 13'sd2964}},
{{7'sd35, 13'sd-3012, 13'sd2849}, {11'sd-822, 12'sd1065, 6'sd21}, {13'sd2617, 13'sd2110, 13'sd3430}},
{{13'sd-2230, 10'sd474, 13'sd2049}, {13'sd-2744, 10'sd509, 13'sd-2686}, {13'sd-2526, 12'sd-1637, 8'sd105}},
{{14'sd-6453, 13'sd-2260, 13'sd-3397}, {12'sd-1512, 12'sd1454, 6'sd18}, {11'sd-602, 14'sd4193, 12'sd1046}},
{{9'sd203, 12'sd1641, 13'sd-2518}, {12'sd-1082, 10'sd437, 9'sd248}, {11'sd598, 12'sd-1405, 12'sd-1034}},
{{12'sd1302, 10'sd408, 13'sd2354}, {13'sd2239, 10'sd-500, 11'sd802}, {12'sd-1919, 12'sd1928, 13'sd2123}},
{{12'sd1930, 13'sd2300, 13'sd-2272}, {13'sd3661, 11'sd-560, 13'sd-3044}, {12'sd1637, 13'sd-2854, 12'sd-1714}},
{{12'sd-1681, 12'sd-2019, 10'sd-325}, {12'sd1247, 12'sd-1209, 13'sd3013}, {13'sd3002, 12'sd-1653, 13'sd2794}},
{{13'sd-2368, 11'sd-724, 13'sd-3539}, {13'sd-2294, 13'sd-3493, 12'sd-1108}, {12'sd-1498, 13'sd-3154, 13'sd-2286}},
{{14'sd6178, 13'sd2105, 11'sd878}, {12'sd1640, 10'sd-453, 12'sd1451}, {11'sd1021, 12'sd-1928, 11'sd990}},
{{13'sd2423, 11'sd860, 12'sd1698}, {12'sd-1239, 9'sd-147, 12'sd1389}, {12'sd1664, 12'sd1746, 11'sd-622}},
{{12'sd1804, 12'sd-1743, 13'sd-2234}, {12'sd1116, 9'sd-146, 11'sd-853}, {12'sd1316, 12'sd1410, 12'sd-1957}},
{{13'sd-2756, 1'sd0, 12'sd-1801}, {8'sd-100, 13'sd-2436, 12'sd-1896}, {9'sd249, 13'sd2659, 13'sd2125}},
{{13'sd2067, 12'sd-2037, 12'sd1965}, {13'sd2114, 12'sd-1891, 12'sd1461}, {12'sd-1940, 12'sd1816, 11'sd-1014}},
{{12'sd1400, 13'sd2382, 13'sd2557}, {10'sd-293, 12'sd1899, 13'sd2268}, {11'sd-1007, 12'sd-1984, 12'sd1328}},
{{13'sd2955, 11'sd-766, 11'sd677}, {12'sd-1130, 12'sd1570, 9'sd225}, {12'sd1139, 12'sd1132, 13'sd-3299}},
{{12'sd1924, 12'sd2037, 13'sd3962}, {12'sd1240, 12'sd1545, 13'sd3900}, {14'sd4650, 12'sd1802, 14'sd5909}},
{{7'sd-59, 12'sd-1124, 12'sd1735}, {12'sd1896, 13'sd2507, 12'sd1315}, {12'sd1449, 11'sd-585, 12'sd1505}},
{{9'sd-196, 12'sd1049, 12'sd-1708}, {11'sd585, 13'sd-2120, 11'sd-926}, {13'sd2271, 12'sd1169, 10'sd-451}},
{{13'sd-3496, 9'sd-242, 13'sd-2464}, {12'sd1057, 11'sd-616, 12'sd-1564}, {12'sd1782, 13'sd-3530, 13'sd-2089}},
{{12'sd1055, 12'sd1487, 11'sd606}, {12'sd-1057, 11'sd557, 12'sd-1533}, {11'sd557, 13'sd2438, 12'sd-1946}},
{{12'sd-1813, 12'sd-1900, 10'sd-475}, {12'sd1727, 13'sd3470, 13'sd2772}, {13'sd2133, 13'sd2866, 8'sd82}},
{{13'sd3203, 12'sd1603, 10'sd506}, {13'sd2907, 12'sd-1952, 13'sd2216}, {13'sd2151, 13'sd2437, 13'sd2856}},
{{14'sd-4541, 13'sd-3570, 12'sd-1220}, {12'sd-1763, 13'sd-3856, 12'sd-1436}, {13'sd-2223, 13'sd-3854, 13'sd-3546}}},
{
{{11'sd863, 12'sd-1963, 12'sd1160}, {12'sd1486, 12'sd-1771, 12'sd-1065}, {11'sd742, 12'sd-1855, 13'sd2170}},
{{11'sd1002, 11'sd-993, 8'sd86}, {13'sd2139, 12'sd-1294, 13'sd2288}, {11'sd-840, 9'sd-243, 10'sd-263}},
{{12'sd-1378, 12'sd2012, 12'sd-2040}, {13'sd2219, 11'sd972, 9'sd238}, {12'sd1256, 11'sd-552, 13'sd2307}},
{{11'sd580, 11'sd-840, 12'sd1908}, {12'sd-1858, 11'sd520, 13'sd-2083}, {12'sd-1448, 12'sd1795, 12'sd-1616}},
{{9'sd-248, 13'sd-2268, 12'sd1513}, {13'sd-2772, 12'sd1820, 12'sd1721}, {12'sd-1951, 10'sd-481, 10'sd327}},
{{13'sd-2332, 9'sd165, 11'sd691}, {12'sd-1515, 13'sd2442, 11'sd645}, {12'sd1585, 12'sd1074, 9'sd-209}},
{{13'sd-2348, 9'sd217, 11'sd669}, {9'sd-225, 12'sd-1378, 10'sd-430}, {12'sd-1636, 13'sd-3136, 12'sd-1528}},
{{11'sd-942, 12'sd1780, 12'sd-1038}, {11'sd-735, 13'sd-2802, 13'sd2255}, {12'sd-1729, 10'sd-357, 13'sd2526}},
{{12'sd-1774, 10'sd-337, 12'sd-1919}, {10'sd-387, 11'sd-533, 9'sd155}, {13'sd2479, 12'sd1100, 10'sd490}},
{{12'sd-1625, 12'sd1123, 12'sd-1719}, {12'sd-1996, 10'sd277, 13'sd2374}, {12'sd1848, 12'sd1421, 13'sd-2485}},
{{12'sd1628, 9'sd-245, 12'sd-1793}, {11'sd764, 10'sd449, 11'sd566}, {12'sd-1967, 13'sd2295, 10'sd391}},
{{12'sd-1310, 13'sd-2629, 13'sd2327}, {12'sd1512, 11'sd978, 7'sd-52}, {13'sd2715, 11'sd-601, 13'sd3108}},
{{13'sd3488, 11'sd-917, 12'sd2007}, {12'sd1765, 13'sd2710, 13'sd2487}, {13'sd2276, 12'sd-1225, 12'sd1785}},
{{12'sd-1627, 12'sd1232, 8'sd86}, {12'sd-1664, 13'sd-2509, 13'sd-2799}, {11'sd969, 12'sd1187, 10'sd463}},
{{13'sd-3636, 9'sd227, 12'sd1216}, {14'sd-4374, 9'sd-230, 12'sd1216}, {12'sd-1890, 14'sd-4783, 13'sd-2795}},
{{10'sd-399, 12'sd2007, 12'sd1413}, {8'sd-87, 10'sd-509, 13'sd3199}, {12'sd1884, 8'sd96, 13'sd3222}},
{{12'sd-1713, 8'sd-73, 12'sd1028}, {11'sd772, 12'sd-1146, 12'sd2022}, {13'sd2554, 12'sd-1617, 13'sd-2300}},
{{12'sd-1647, 13'sd-2963, 11'sd673}, {11'sd-566, 11'sd-529, 13'sd2476}, {12'sd1420, 6'sd25, 10'sd441}},
{{11'sd-959, 12'sd1452, 13'sd-2453}, {12'sd-1597, 11'sd-962, 12'sd-1031}, {13'sd-2724, 12'sd-1662, 10'sd-358}},
{{11'sd585, 7'sd55, 9'sd176}, {12'sd1826, 12'sd-1723, 13'sd2328}, {12'sd-1943, 11'sd840, 9'sd178}},
{{13'sd-2375, 13'sd2395, 10'sd493}, {11'sd-959, 12'sd-1548, 12'sd-1448}, {11'sd771, 13'sd2139, 13'sd-2374}},
{{12'sd1406, 12'sd1850, 12'sd1092}, {4'sd-5, 12'sd1690, 11'sd965}, {12'sd-1565, 12'sd-1572, 12'sd-1031}},
{{13'sd2721, 13'sd2973, 11'sd-891}, {10'sd336, 12'sd1193, 13'sd2130}, {12'sd-1962, 12'sd-1576, 9'sd168}},
{{13'sd-2121, 12'sd-2024, 12'sd-1083}, {13'sd-2327, 11'sd-911, 10'sd-281}, {12'sd1205, 12'sd-1247, 12'sd-1080}},
{{12'sd1575, 12'sd-1115, 13'sd2124}, {11'sd896, 12'sd-1834, 12'sd1137}, {12'sd-1077, 12'sd1197, 13'sd-2159}},
{{11'sd-918, 12'sd-1184, 13'sd-2189}, {12'sd-1111, 12'sd-1838, 12'sd1035}, {12'sd1861, 12'sd1177, 13'sd2786}},
{{11'sd660, 12'sd-1602, 12'sd-1994}, {13'sd3190, 11'sd-521, 13'sd-2266}, {13'sd3483, 11'sd947, 12'sd1075}},
{{4'sd6, 13'sd-2152, 11'sd887}, {9'sd188, 12'sd-1077, 11'sd900}, {13'sd-3326, 13'sd-2877, 7'sd-61}},
{{12'sd1310, 12'sd-1847, 12'sd-2016}, {12'sd1563, 13'sd-2285, 13'sd-2543}, {10'sd-438, 11'sd562, 13'sd-2907}},
{{9'sd213, 12'sd-1507, 12'sd-2031}, {11'sd-710, 12'sd1854, 13'sd-3063}, {10'sd-499, 7'sd-38, 13'sd-2840}},
{{10'sd350, 10'sd-287, 11'sd-590}, {13'sd2224, 12'sd1611, 9'sd-167}, {13'sd2471, 12'sd-1154, 13'sd-2370}},
{{12'sd-1800, 11'sd-943, 13'sd2479}, {11'sd1021, 4'sd6, 12'sd-1856}, {12'sd-1663, 8'sd77, 12'sd-1663}},
{{10'sd-419, 13'sd2124, 9'sd-234}, {12'sd1531, 12'sd1993, 13'sd-2808}, {7'sd56, 13'sd2544, 13'sd2245}},
{{12'sd-1348, 11'sd597, 10'sd-445}, {12'sd1864, 11'sd-602, 10'sd349}, {12'sd1332, 9'sd250, 10'sd428}},
{{10'sd427, 11'sd615, 13'sd-2568}, {13'sd-2255, 11'sd935, 10'sd-361}, {9'sd143, 13'sd-2224, 13'sd-2413}},
{{12'sd-1424, 12'sd-1202, 11'sd982}, {12'sd1554, 8'sd-98, 12'sd-1280}, {11'sd867, 12'sd-1295, 10'sd-280}},
{{13'sd3577, 10'sd-488, 12'sd-1102}, {11'sd665, 11'sd-655, 11'sd908}, {12'sd-1321, 11'sd1005, 9'sd-215}},
{{12'sd1769, 10'sd350, 12'sd1256}, {12'sd1270, 12'sd-1917, 12'sd1523}, {12'sd1367, 12'sd2038, 8'sd70}},
{{12'sd1105, 12'sd1728, 13'sd2401}, {12'sd1107, 12'sd-1425, 13'sd-2269}, {13'sd-2577, 10'sd-464, 11'sd-677}},
{{11'sd-957, 13'sd2791, 11'sd-904}, {12'sd-1626, 7'sd-45, 11'sd778}, {12'sd-1086, 12'sd2027, 12'sd-1145}},
{{12'sd-1902, 13'sd-2509, 10'sd-465}, {11'sd650, 13'sd-2102, 12'sd-1390}, {12'sd1777, 12'sd2017, 11'sd-938}},
{{13'sd2780, 13'sd2219, 12'sd1317}, {12'sd-1068, 6'sd-28, 10'sd-353}, {13'sd2672, 13'sd4071, 12'sd-1577}},
{{8'sd97, 12'sd-1523, 11'sd738}, {9'sd-219, 12'sd-1712, 13'sd-3622}, {12'sd-1084, 12'sd1773, 12'sd-1538}},
{{10'sd-341, 9'sd254, 12'sd1211}, {14'sd5358, 13'sd2427, 12'sd-1257}, {14'sd7890, 13'sd3800, 14'sd5525}},
{{12'sd-1142, 8'sd-100, 13'sd-2566}, {13'sd-2094, 12'sd1989, 13'sd-2113}, {11'sd-715, 11'sd568, 12'sd1863}},
{{11'sd945, 13'sd2810, 12'sd1851}, {13'sd2087, 8'sd-90, 12'sd-1968}, {12'sd1726, 12'sd-1269, 13'sd2765}},
{{13'sd2207, 9'sd188, 11'sd-991}, {12'sd-1125, 13'sd2228, 12'sd1906}, {12'sd1401, 13'sd2526, 9'sd-204}},
{{13'sd-2188, 12'sd-1848, 10'sd336}, {12'sd-1388, 12'sd1759, 12'sd-1575}, {13'sd-3625, 10'sd-327, 11'sd-542}},
{{13'sd-3882, 13'sd-2199, 11'sd-706}, {13'sd-3732, 13'sd-2279, 11'sd821}, {12'sd-1490, 12'sd1251, 12'sd2044}},
{{13'sd2618, 12'sd1082, 12'sd-1651}, {10'sd462, 9'sd-204, 13'sd2684}, {12'sd1429, 13'sd2054, 10'sd-466}},
{{5'sd10, 11'sd941, 12'sd-1722}, {12'sd1541, 12'sd1978, 7'sd-35}, {11'sd640, 11'sd981, 9'sd-163}},
{{11'sd764, 13'sd2488, 9'sd-149}, {12'sd1621, 10'sd271, 11'sd787}, {13'sd2415, 12'sd-1535, 8'sd90}},
{{13'sd2119, 11'sd-685, 11'sd-750}, {11'sd733, 11'sd806, 13'sd-2443}, {12'sd1438, 12'sd-1869, 9'sd216}},
{{8'sd-81, 11'sd-861, 7'sd51}, {12'sd1908, 13'sd2329, 11'sd-524}, {11'sd579, 11'sd-927, 13'sd2633}},
{{13'sd3161, 12'sd1337, 9'sd-245}, {11'sd-1001, 12'sd-1881, 12'sd-1079}, {5'sd8, 12'sd-1273, 10'sd511}},
{{13'sd3323, 12'sd-1271, 10'sd380}, {11'sd778, 13'sd2354, 13'sd2307}, {11'sd-673, 10'sd-407, 12'sd-1293}},
{{11'sd-524, 11'sd546, 11'sd772}, {12'sd-1055, 12'sd-1803, 12'sd-1181}, {11'sd-705, 11'sd959, 9'sd182}},
{{11'sd967, 10'sd-486, 11'sd-771}, {7'sd45, 12'sd-1068, 13'sd2257}, {13'sd-2444, 12'sd1586, 12'sd1759}},
{{13'sd2245, 13'sd-2723, 12'sd-1284}, {12'sd1453, 10'sd342, 10'sd-495}, {13'sd2166, 13'sd2179, 12'sd-1421}},
{{5'sd-8, 12'sd1499, 6'sd22}, {12'sd-2001, 12'sd1349, 13'sd-2332}, {9'sd-179, 12'sd1406, 13'sd3048}},
{{11'sd-710, 13'sd2169, 12'sd1098}, {12'sd2043, 12'sd-1062, 9'sd224}, {9'sd-160, 12'sd-1811, 12'sd-1152}},
{{11'sd-606, 13'sd2205, 12'sd-1047}, {12'sd1293, 12'sd-1849, 12'sd-1620}, {12'sd-1130, 13'sd2824, 10'sd294}},
{{12'sd2036, 13'sd2707, 11'sd752}, {11'sd-864, 12'sd-1316, 12'sd-1723}, {10'sd-292, 12'sd-1677, 12'sd-1461}},
{{13'sd2250, 13'sd-2326, 12'sd-1865}, {12'sd-1812, 12'sd-1595, 13'sd-2969}, {13'sd-2380, 13'sd-3508, 12'sd-1029}}},
{
{{13'sd-2181, 9'sd-204, 12'sd1703}, {12'sd1068, 12'sd1821, 12'sd1562}, {12'sd-1497, 12'sd1593, 12'sd-1240}},
{{12'sd-1317, 11'sd901, 5'sd8}, {11'sd-869, 10'sd483, 12'sd1569}, {12'sd-1181, 12'sd-1302, 12'sd1355}},
{{12'sd1090, 13'sd-2423, 11'sd739}, {13'sd2757, 13'sd2203, 12'sd-1928}, {11'sd-644, 8'sd95, 12'sd-1817}},
{{12'sd1947, 13'sd-2135, 13'sd2423}, {9'sd-215, 8'sd97, 12'sd-1208}, {12'sd1460, 11'sd-627, 11'sd-564}},
{{14'sd4126, 13'sd2995, 13'sd2981}, {12'sd1632, 11'sd-1018, 11'sd-609}, {13'sd3256, 13'sd2520, 12'sd-1891}},
{{13'sd-3427, 4'sd-7, 13'sd2999}, {10'sd-310, 11'sd906, 13'sd2498}, {12'sd1840, 11'sd-721, 6'sd23}},
{{12'sd1473, 11'sd-831, 13'sd3889}, {10'sd-392, 12'sd-1248, 13'sd-3496}, {12'sd1544, 14'sd-4636, 14'sd-4273}},
{{12'sd-1492, 11'sd-939, 12'sd1895}, {12'sd-1541, 11'sd889, 11'sd-813}, {13'sd2547, 11'sd-992, 13'sd2099}},
{{13'sd-2885, 13'sd-2954, 11'sd-921}, {12'sd1816, 11'sd-559, 10'sd487}, {12'sd-1761, 12'sd-1190, 10'sd391}},
{{13'sd2555, 12'sd1703, 9'sd217}, {11'sd-764, 13'sd-2137, 12'sd-1809}, {13'sd3591, 13'sd-2713, 9'sd138}},
{{11'sd-572, 13'sd2717, 12'sd1725}, {9'sd242, 10'sd496, 12'sd1731}, {11'sd-694, 10'sd-395, 13'sd2472}},
{{12'sd-1693, 13'sd2560, 2'sd1}, {9'sd193, 13'sd2876, 10'sd-266}, {12'sd1168, 13'sd2076, 12'sd-1290}},
{{13'sd3127, 12'sd1964, 9'sd212}, {12'sd1713, 13'sd-2419, 12'sd-2001}, {12'sd-1493, 12'sd1628, 9'sd190}},
{{13'sd2798, 10'sd416, 13'sd2635}, {13'sd-2262, 11'sd-681, 9'sd233}, {12'sd-2041, 12'sd1505, 13'sd-2469}},
{{13'sd3516, 12'sd2016, 13'sd3175}, {12'sd1123, 11'sd552, 13'sd-3056}, {13'sd3186, 13'sd3974, 12'sd-1037}},
{{12'sd1273, 13'sd-2736, 11'sd612}, {13'sd-2327, 13'sd-2708, 11'sd-574}, {11'sd-682, 12'sd1469, 13'sd-2977}},
{{13'sd2628, 13'sd-2140, 13'sd3074}, {13'sd2366, 11'sd-623, 12'sd-1703}, {12'sd1910, 12'sd-1689, 13'sd2607}},
{{6'sd-21, 12'sd-1337, 12'sd1517}, {11'sd-705, 12'sd-1088, 9'sd-135}, {13'sd-2854, 13'sd-3678, 12'sd-1612}},
{{11'sd-945, 13'sd2143, 13'sd-2211}, {12'sd1280, 11'sd834, 11'sd953}, {10'sd-321, 11'sd1020, 12'sd-1565}},
{{7'sd-63, 13'sd-2409, 13'sd2304}, {9'sd227, 12'sd-1421, 13'sd2603}, {13'sd-2815, 11'sd-694, 13'sd-2650}},
{{12'sd1256, 13'sd2674, 13'sd3207}, {12'sd1637, 12'sd1928, 12'sd1080}, {12'sd-2026, 12'sd-1215, 13'sd2625}},
{{11'sd942, 13'sd2404, 13'sd3168}, {11'sd-860, 13'sd2195, 12'sd-1107}, {11'sd647, 12'sd-2017, 12'sd1140}},
{{11'sd1002, 12'sd-1866, 13'sd2786}, {13'sd2873, 13'sd-2831, 12'sd1435}, {9'sd-216, 12'sd-1612, 12'sd1911}},
{{12'sd1174, 12'sd-1131, 13'sd2975}, {9'sd-241, 11'sd-659, 13'sd2491}, {11'sd963, 9'sd-252, 9'sd153}},
{{11'sd-964, 12'sd-1216, 12'sd1220}, {13'sd2724, 11'sd686, 12'sd-2010}, {12'sd-1479, 13'sd-3165, 11'sd-781}},
{{12'sd1808, 12'sd1205, 10'sd258}, {11'sd825, 9'sd-183, 12'sd-1116}, {12'sd1550, 12'sd-1369, 10'sd-423}},
{{13'sd-2527, 13'sd-2925, 13'sd-2950}, {10'sd-367, 11'sd933, 11'sd-893}, {13'sd-2489, 11'sd-604, 11'sd980}},
{{13'sd-2187, 12'sd1128, 12'sd-1612}, {10'sd335, 13'sd2555, 12'sd-1328}, {4'sd5, 12'sd1398, 11'sd-959}},
{{13'sd3777, 11'sd867, 13'sd-2170}, {12'sd1689, 13'sd2164, 11'sd758}, {9'sd194, 11'sd523, 12'sd1894}},
{{13'sd-3222, 13'sd-2498, 11'sd705}, {13'sd-3377, 12'sd1231, 10'sd396}, {11'sd-954, 13'sd2917, 13'sd2634}},
{{12'sd-1349, 11'sd-873, 12'sd1254}, {11'sd605, 12'sd1193, 6'sd-26}, {8'sd-72, 13'sd-2681, 13'sd2739}},
{{12'sd1128, 8'sd96, 13'sd2148}, {13'sd2659, 11'sd891, 12'sd-1736}, {12'sd1452, 12'sd-2024, 7'sd47}},
{{12'sd-1899, 11'sd657, 11'sd1007}, {11'sd-580, 12'sd1984, 11'sd734}, {10'sd-360, 13'sd-2234, 12'sd-1441}},
{{13'sd-2454, 12'sd-1110, 10'sd466}, {11'sd-705, 13'sd2668, 12'sd1712}, {10'sd349, 13'sd2574, 11'sd-856}},
{{9'sd142, 12'sd1064, 13'sd-2158}, {11'sd-877, 10'sd282, 12'sd1673}, {12'sd-1757, 13'sd-2440, 13'sd2987}},
{{13'sd-2353, 9'sd130, 9'sd-213}, {11'sd-572, 13'sd-2997, 11'sd-917}, {11'sd-999, 12'sd-1415, 13'sd-2274}},
{{9'sd-231, 12'sd-1337, 11'sd661}, {13'sd-2394, 13'sd-2440, 13'sd2859}, {13'sd-3699, 11'sd-1023, 10'sd337}},
{{7'sd-49, 10'sd-409, 12'sd-1595}, {12'sd-1345, 11'sd-731, 10'sd393}, {13'sd-2837, 12'sd-1178, 12'sd-1702}},
{{12'sd-1412, 12'sd1229, 11'sd-864}, {12'sd1248, 12'sd-1774, 13'sd2759}, {12'sd-1614, 13'sd-2288, 12'sd-1714}},
{{12'sd-1039, 13'sd-2151, 12'sd-1854}, {10'sd502, 12'sd1252, 12'sd-1277}, {13'sd2924, 12'sd-1764, 7'sd-45}},
{{12'sd-1173, 13'sd-3335, 7'sd-33}, {12'sd-1932, 12'sd-1310, 12'sd-1765}, {11'sd-728, 13'sd-3093, 13'sd-2655}},
{{12'sd1573, 11'sd719, 12'sd1776}, {11'sd873, 12'sd-1216, 11'sd645}, {12'sd-1435, 12'sd1097, 13'sd-2949}},
{{12'sd1481, 13'sd3221, 13'sd-2121}, {10'sd457, 9'sd-240, 12'sd1772}, {13'sd-2375, 13'sd2786, 11'sd-935}},
{{15'sd9733, 11'sd623, 14'sd5124}, {12'sd-1359, 14'sd-4601, 11'sd-735}, {13'sd2517, 12'sd-1870, 13'sd2721}},
{{13'sd2054, 13'sd-2958, 7'sd47}, {10'sd410, 11'sd801, 10'sd346}, {12'sd1835, 12'sd-1208, 12'sd1347}},
{{13'sd2348, 10'sd-336, 12'sd1390}, {12'sd-1878, 12'sd-1578, 13'sd2980}, {13'sd-2439, 12'sd1190, 9'sd134}},
{{13'sd-3643, 13'sd-3038, 11'sd705}, {8'sd66, 12'sd1267, 12'sd-1093}, {13'sd-3252, 10'sd-436, 11'sd814}},
{{12'sd-1149, 13'sd3403, 12'sd1574}, {13'sd-2785, 12'sd-1715, 13'sd-2477}, {13'sd-2850, 10'sd-283, 12'sd1151}},
{{13'sd-3366, 11'sd-932, 10'sd267}, {13'sd-3192, 10'sd-509, 13'sd2709}, {12'sd-1602, 12'sd-1981, 12'sd1191}},
{{13'sd-3082, 10'sd320, 11'sd-833}, {13'sd-3659, 12'sd1271, 13'sd3640}, {7'sd-58, 13'sd2127, 13'sd3006}},
{{8'sd-118, 13'sd3272, 12'sd-1705}, {12'sd-1513, 9'sd-147, 8'sd-71}, {7'sd-38, 11'sd683, 13'sd-2472}},
{{10'sd-346, 7'sd34, 10'sd-442}, {10'sd437, 13'sd2222, 12'sd-1311}, {11'sd-942, 9'sd-249, 11'sd-706}},
{{11'sd-864, 12'sd1093, 13'sd-2153}, {13'sd3365, 11'sd-586, 13'sd-2546}, {13'sd3656, 13'sd3266, 13'sd-2613}},
{{13'sd2664, 9'sd-253, 13'sd2811}, {12'sd-2002, 13'sd2353, 13'sd2536}, {11'sd823, 10'sd-444, 12'sd1374}},
{{10'sd-405, 13'sd3144, 10'sd-403}, {12'sd-1355, 10'sd-394, 13'sd-3936}, {13'sd-3281, 11'sd-729, 6'sd23}},
{{12'sd1126, 13'sd-2593, 10'sd311}, {11'sd-975, 11'sd526, 13'sd2504}, {9'sd212, 10'sd388, 13'sd3082}},
{{14'sd5101, 12'sd1287, 7'sd-51}, {13'sd-3107, 13'sd3528, 13'sd-2783}, {14'sd4148, 12'sd1991, 13'sd-2768}},
{{7'sd61, 13'sd-3172, 11'sd767}, {13'sd2464, 12'sd-1610, 13'sd-3391}, {11'sd708, 13'sd-3053, 13'sd-2645}},
{{12'sd-1601, 12'sd1220, 12'sd2038}, {10'sd-350, 9'sd-134, 12'sd-1890}, {12'sd1256, 11'sd517, 12'sd1627}},
{{13'sd-3458, 12'sd-1743, 10'sd263}, {11'sd-927, 12'sd1615, 11'sd868}, {15'sd-8405, 12'sd-1499, 12'sd-1643}},
{{12'sd-1943, 10'sd424, 12'sd-1543}, {10'sd-360, 12'sd-1121, 12'sd1552}, {12'sd1587, 11'sd-906, 11'sd-651}},
{{12'sd-1752, 12'sd-2006, 13'sd-3106}, {13'sd2383, 13'sd2206, 12'sd1968}, {11'sd-791, 11'sd-889, 13'sd-2263}},
{{8'sd-66, 12'sd-1350, 13'sd2261}, {9'sd-222, 13'sd-2287, 10'sd-267}, {10'sd-478, 13'sd-3161, 12'sd-1040}},
{{13'sd3591, 11'sd-957, 13'sd3402}, {11'sd-999, 12'sd1699, 13'sd3077}, {12'sd1470, 13'sd2234, 11'sd-747}}},
{
{{13'sd2140, 12'sd-1741, 8'sd120}, {9'sd244, 12'sd1489, 13'sd-2657}, {12'sd-1985, 12'sd-1634, 10'sd-411}},
{{10'sd-326, 13'sd2186, 11'sd-831}, {12'sd-1507, 11'sd698, 11'sd761}, {10'sd497, 12'sd-1417, 12'sd1045}},
{{12'sd-1748, 10'sd-448, 11'sd693}, {13'sd-2378, 13'sd2531, 13'sd2195}, {11'sd-594, 12'sd1462, 13'sd2354}},
{{13'sd2116, 11'sd983, 12'sd1117}, {13'sd2854, 13'sd2798, 12'sd-1351}, {11'sd935, 13'sd2901, 12'sd-1335}},
{{13'sd2866, 13'sd3984, 12'sd2013}, {11'sd-644, 13'sd2737, 12'sd-1262}, {14'sd4181, 14'sd4696, 12'sd1438}},
{{13'sd2180, 10'sd503, 12'sd-1192}, {10'sd405, 9'sd-198, 12'sd1674}, {11'sd-704, 12'sd1176, 13'sd-2752}},
{{12'sd1330, 13'sd3787, 13'sd2522}, {13'sd2576, 11'sd543, 13'sd2898}, {13'sd2957, 12'sd-1362, 11'sd-595}},
{{12'sd1820, 13'sd2551, 11'sd-794}, {13'sd-2205, 12'sd1062, 13'sd-2578}, {13'sd-2518, 11'sd-815, 12'sd1493}},
{{11'sd823, 12'sd1585, 11'sd-782}, {11'sd-581, 12'sd-1178, 12'sd1711}, {12'sd-1216, 10'sd-481, 12'sd1126}},
{{12'sd-1912, 12'sd1162, 12'sd1264}, {13'sd-2484, 12'sd-1356, 13'sd2774}, {13'sd2196, 11'sd742, 12'sd1715}},
{{10'sd-266, 13'sd2356, 10'sd367}, {8'sd71, 11'sd-995, 12'sd1717}, {12'sd2018, 12'sd1387, 10'sd432}},
{{11'sd-844, 12'sd-2036, 13'sd-2310}, {9'sd197, 10'sd470, 10'sd-381}, {10'sd367, 11'sd599, 10'sd-468}},
{{11'sd-581, 12'sd1402, 12'sd1640}, {13'sd2863, 13'sd3670, 13'sd2675}, {10'sd509, 10'sd307, 8'sd70}},
{{12'sd-1947, 11'sd-664, 11'sd558}, {13'sd-2291, 11'sd-923, 12'sd-1113}, {11'sd986, 13'sd2308, 11'sd612}},
{{10'sd-419, 12'sd1576, 10'sd-375}, {12'sd-1585, 12'sd-1324, 11'sd-529}, {11'sd-674, 11'sd-794, 14'sd4994}},
{{13'sd2833, 12'sd1710, 12'sd1158}, {10'sd-328, 13'sd-2133, 12'sd-1476}, {13'sd-2699, 12'sd-1070, 12'sd-1071}},
{{11'sd531, 12'sd2015, 12'sd1122}, {12'sd-1484, 13'sd-2869, 11'sd-932}, {12'sd1430, 10'sd427, 12'sd-1455}},
{{12'sd-1252, 11'sd833, 12'sd1213}, {13'sd2631, 12'sd1553, 13'sd3269}, {12'sd1565, 13'sd3451, 12'sd2008}},
{{13'sd-2172, 11'sd-785, 10'sd330}, {13'sd2551, 12'sd-1656, 12'sd-1684}, {13'sd2119, 12'sd1748, 10'sd398}},
{{12'sd-1649, 12'sd1731, 12'sd1072}, {8'sd83, 11'sd950, 10'sd-302}, {13'sd-2854, 10'sd388, 10'sd434}},
{{12'sd1178, 13'sd2099, 13'sd-2800}, {11'sd-822, 12'sd-1569, 12'sd-1791}, {11'sd-990, 12'sd1346, 13'sd2404}},
{{12'sd-1333, 10'sd-494, 10'sd-324}, {11'sd-1020, 12'sd-1596, 11'sd-881}, {11'sd-744, 11'sd515, 12'sd1696}},
{{7'sd55, 10'sd-380, 13'sd2603}, {12'sd-1494, 12'sd-1877, 11'sd586}, {11'sd-955, 11'sd-792, 12'sd-1117}},
{{13'sd2105, 11'sd529, 12'sd-1932}, {13'sd-2054, 10'sd382, 11'sd996}, {12'sd-1559, 11'sd844, 12'sd1420}},
{{12'sd-1083, 12'sd-1662, 12'sd-1814}, {12'sd-1765, 13'sd2366, 13'sd-2247}, {12'sd1286, 5'sd13, 12'sd-1617}},
{{12'sd1210, 13'sd2232, 13'sd2881}, {13'sd-2330, 12'sd-1500, 12'sd1734}, {12'sd1561, 13'sd2255, 11'sd-635}},
{{11'sd-660, 11'sd689, 13'sd2354}, {7'sd-62, 12'sd1446, 13'sd2208}, {13'sd4081, 11'sd1015, 11'sd-700}},
{{11'sd-908, 11'sd860, 11'sd936}, {13'sd2733, 13'sd2470, 11'sd972}, {11'sd-829, 13'sd2814, 12'sd1214}},
{{12'sd1738, 10'sd425, 11'sd812}, {13'sd-2477, 12'sd-1676, 10'sd-289}, {12'sd-1246, 11'sd-553, 12'sd1129}},
{{11'sd-574, 12'sd-1892, 9'sd159}, {11'sd-1001, 11'sd626, 10'sd350}, {12'sd1276, 11'sd-624, 12'sd-1771}},
{{12'sd-1587, 12'sd-1205, 12'sd-1913}, {9'sd-154, 13'sd-2233, 13'sd-2365}, {13'sd-2726, 12'sd1303, 12'sd1394}},
{{11'sd-698, 11'sd-805, 3'sd-3}, {13'sd-2876, 11'sd-626, 12'sd-1641}, {12'sd-1738, 9'sd239, 12'sd-1817}},
{{11'sd551, 12'sd-1599, 10'sd-285}, {12'sd1735, 12'sd-2028, 11'sd866}, {11'sd861, 10'sd425, 11'sd-912}},
{{11'sd-889, 11'sd810, 12'sd1111}, {10'sd428, 9'sd145, 12'sd-1740}, {13'sd-2260, 7'sd-62, 12'sd-1243}},
{{10'sd-404, 13'sd-2116, 12'sd-1220}, {12'sd1973, 12'sd1665, 13'sd-3410}, {10'sd322, 13'sd-2652, 12'sd1659}},
{{12'sd-1265, 12'sd-1393, 11'sd-768}, {13'sd-2496, 11'sd1023, 13'sd-2970}, {13'sd-2346, 11'sd977, 13'sd2367}},
{{12'sd1436, 12'sd-1488, 12'sd-1104}, {12'sd1266, 12'sd-1931, 11'sd-724}, {12'sd1347, 14'sd-4168, 11'sd907}},
{{11'sd-551, 11'sd941, 12'sd1132}, {12'sd1031, 13'sd2615, 13'sd2668}, {12'sd1741, 13'sd2832, 13'sd3145}},
{{11'sd865, 11'sd749, 9'sd219}, {9'sd-167, 10'sd275, 12'sd-1038}, {7'sd-52, 12'sd1923, 13'sd-2320}},
{{10'sd391, 12'sd1463, 13'sd2198}, {12'sd2044, 13'sd-2462, 9'sd148}, {12'sd1170, 12'sd1148, 9'sd-158}},
{{11'sd-625, 12'sd-1472, 10'sd258}, {12'sd1507, 10'sd-260, 12'sd-1526}, {12'sd-1661, 13'sd3350, 12'sd-1242}},
{{13'sd2082, 13'sd-2498, 13'sd2324}, {11'sd-544, 13'sd2878, 12'sd1040}, {7'sd-35, 13'sd2253, 12'sd1052}},
{{11'sd-847, 13'sd2053, 13'sd3656}, {12'sd-1475, 13'sd2556, 10'sd486}, {10'sd-401, 12'sd1500, 8'sd-98}},
{{11'sd843, 10'sd-477, 7'sd44}, {13'sd2988, 12'sd1744, 10'sd-296}, {13'sd2499, 13'sd3139, 12'sd1465}},
{{12'sd1027, 12'sd1120, 12'sd-1832}, {12'sd1885, 13'sd2420, 12'sd1617}, {13'sd2540, 12'sd1805, 12'sd1309}},
{{13'sd-2627, 13'sd2266, 13'sd-2454}, {13'sd-2502, 11'sd-802, 13'sd2222}, {10'sd-290, 13'sd2562, 11'sd-1006}},
{{13'sd3195, 12'sd-1501, 11'sd964}, {12'sd1880, 13'sd-2106, 11'sd705}, {11'sd-957, 12'sd-1605, 12'sd-1990}},
{{12'sd-1340, 12'sd-1587, 12'sd1835}, {12'sd1227, 12'sd1643, 6'sd-16}, {11'sd947, 12'sd1369, 12'sd1329}},
{{11'sd754, 12'sd-1113, 12'sd1863}, {13'sd2601, 11'sd-865, 11'sd-846}, {12'sd1988, 10'sd374, 13'sd-2561}},
{{12'sd2026, 12'sd-1093, 13'sd2370}, {12'sd-1369, 11'sd-927, 7'sd-43}, {12'sd1049, 12'sd-1720, 12'sd-1330}},
{{11'sd907, 12'sd-1528, 13'sd-2095}, {13'sd-2841, 12'sd1446, 13'sd2636}, {8'sd83, 13'sd-2387, 10'sd422}},
{{12'sd1647, 13'sd-2552, 12'sd-1680}, {13'sd-2079, 8'sd78, 12'sd1603}, {13'sd-2564, 13'sd-2226, 12'sd-1973}},
{{13'sd-2358, 11'sd617, 11'sd884}, {12'sd1119, 12'sd1422, 12'sd-1298}, {11'sd-797, 11'sd-522, 9'sd-197}},
{{12'sd1413, 13'sd2117, 13'sd-2085}, {9'sd209, 11'sd565, 12'sd1513}, {11'sd754, 8'sd75, 10'sd-483}},
{{11'sd840, 13'sd3085, 13'sd3951}, {13'sd2129, 10'sd-355, 13'sd2294}, {13'sd3042, 10'sd323, 13'sd3714}},
{{11'sd953, 11'sd703, 12'sd-1417}, {13'sd-2445, 12'sd-1998, 13'sd-2797}, {13'sd2236, 12'sd1346, 11'sd963}},
{{13'sd2131, 13'sd2521, 8'sd-91}, {12'sd-1396, 13'sd2215, 13'sd3260}, {11'sd647, 13'sd3792, 13'sd3710}},
{{12'sd1137, 12'sd1223, 11'sd822}, {12'sd1826, 12'sd1303, 10'sd316}, {13'sd2344, 11'sd676, 12'sd-1863}},
{{13'sd-2134, 11'sd-527, 13'sd2071}, {12'sd1125, 12'sd1403, 9'sd176}, {12'sd-1913, 12'sd1030, 12'sd-1927}},
{{12'sd-1062, 12'sd1894, 10'sd-344}, {11'sd794, 11'sd-750, 13'sd3074}, {12'sd-1228, 7'sd-38, 13'sd2550}},
{{13'sd-2417, 13'sd2440, 13'sd-2816}, {12'sd1584, 10'sd303, 12'sd-1292}, {12'sd-1981, 11'sd-848, 8'sd-111}},
{{12'sd-1251, 10'sd289, 12'sd1353}, {12'sd-1748, 12'sd1801, 13'sd2539}, {9'sd152, 12'sd1135, 12'sd1398}},
{{12'sd-1711, 13'sd-2696, 13'sd-3115}, {9'sd-204, 11'sd-637, 12'sd1031}, {10'sd482, 13'sd2242, 8'sd67}},
{{11'sd-568, 13'sd-2670, 12'sd-1655}, {11'sd-927, 12'sd1846, 13'sd-2333}, {12'sd-1747, 13'sd-2776, 13'sd-2833}}},
{
{{11'sd-742, 11'sd-577, 12'sd1971}, {11'sd-547, 12'sd-1288, 12'sd-1698}, {12'sd-1946, 13'sd-2552, 12'sd-1419}},
{{12'sd1041, 11'sd769, 7'sd58}, {12'sd2041, 11'sd602, 12'sd1359}, {11'sd888, 12'sd1427, 13'sd3085}},
{{10'sd-467, 12'sd1927, 13'sd-2504}, {9'sd-217, 12'sd-1779, 13'sd2504}, {11'sd779, 9'sd-218, 12'sd2020}},
{{11'sd785, 12'sd-1709, 12'sd1118}, {13'sd-2525, 11'sd781, 12'sd1832}, {13'sd-2610, 11'sd-819, 13'sd-2790}},
{{11'sd-930, 11'sd753, 13'sd2649}, {11'sd-611, 12'sd1283, 13'sd-2191}, {13'sd-3040, 13'sd-2677, 11'sd513}},
{{12'sd-1222, 13'sd2073, 11'sd-836}, {13'sd-2457, 13'sd3782, 13'sd2209}, {13'sd3482, 12'sd-1328, 11'sd861}},
{{13'sd-3631, 11'sd963, 13'sd2230}, {11'sd-947, 12'sd1060, 12'sd-1488}, {13'sd-3173, 12'sd-1477, 11'sd832}},
{{12'sd1912, 11'sd1011, 11'sd594}, {11'sd-994, 10'sd344, 12'sd1823}, {11'sd-631, 13'sd2145, 11'sd-634}},
{{10'sd-263, 11'sd-566, 13'sd2647}, {13'sd2382, 11'sd672, 10'sd-264}, {11'sd952, 12'sd1435, 13'sd2113}},
{{8'sd127, 10'sd480, 12'sd1746}, {12'sd-1869, 10'sd-277, 7'sd-43}, {12'sd1395, 11'sd871, 13'sd2315}},
{{13'sd-2112, 13'sd-2845, 13'sd2362}, {12'sd-1955, 13'sd-2565, 12'sd1144}, {11'sd-543, 11'sd838, 11'sd1016}},
{{13'sd-2359, 9'sd255, 12'sd-1910}, {11'sd-984, 10'sd343, 13'sd2567}, {9'sd-223, 12'sd-1501, 12'sd1316}},
{{11'sd531, 12'sd1150, 11'sd808}, {13'sd2202, 12'sd-1429, 11'sd715}, {13'sd2341, 12'sd-1138, 13'sd2116}},
{{11'sd-665, 13'sd2383, 12'sd-1054}, {12'sd1929, 12'sd1966, 13'sd2171}, {12'sd-1997, 12'sd1718, 12'sd-1928}},
{{14'sd-4235, 11'sd-586, 11'sd-669}, {13'sd-2361, 13'sd-3463, 13'sd-2096}, {14'sd-5578, 12'sd-2017, 12'sd-1423}},
{{12'sd1470, 11'sd591, 11'sd544}, {12'sd-1429, 11'sd592, 13'sd3051}, {10'sd458, 9'sd199, 13'sd2948}},
{{11'sd763, 9'sd-227, 12'sd-1276}, {10'sd344, 12'sd1212, 11'sd-654}, {12'sd1491, 12'sd1101, 11'sd-782}},
{{13'sd-2225, 11'sd832, 13'sd2570}, {8'sd-83, 12'sd1376, 13'sd3298}, {12'sd-1744, 10'sd444, 11'sd-932}},
{{12'sd1284, 7'sd59, 11'sd757}, {12'sd1796, 12'sd1441, 7'sd35}, {12'sd-1275, 12'sd-1795, 12'sd-1292}},
{{11'sd-985, 11'sd-576, 12'sd-1986}, {12'sd1731, 13'sd2530, 13'sd-2155}, {12'sd-1435, 13'sd-2600, 12'sd-1848}},
{{12'sd-1495, 12'sd1089, 12'sd1031}, {13'sd-2561, 11'sd-884, 12'sd-1093}, {13'sd-2553, 11'sd759, 13'sd-3192}},
{{13'sd2741, 11'sd-704, 11'sd-974}, {13'sd2143, 13'sd2703, 12'sd-1972}, {12'sd2009, 10'sd-390, 10'sd416}},
{{11'sd782, 11'sd785, 12'sd-1695}, {13'sd3153, 12'sd-1071, 11'sd-662}, {11'sd809, 12'sd-1534, 12'sd1124}},
{{12'sd1275, 10'sd316, 12'sd-1754}, {13'sd2645, 12'sd-1749, 12'sd-1839}, {12'sd1905, 12'sd-1740, 11'sd-640}},
{{13'sd2702, 13'sd2112, 11'sd921}, {13'sd2183, 12'sd-1738, 10'sd400}, {13'sd2426, 13'sd2610, 12'sd-1300}},
{{12'sd1828, 13'sd-2640, 11'sd664}, {12'sd1492, 13'sd2255, 10'sd-316}, {13'sd-2209, 11'sd768, 13'sd2404}},
{{14'sd-4353, 13'sd-2411, 11'sd717}, {11'sd741, 9'sd155, 11'sd823}, {13'sd2561, 13'sd2455, 13'sd3315}},
{{10'sd472, 11'sd814, 12'sd1930}, {12'sd-1431, 12'sd-1457, 12'sd-1866}, {13'sd-2880, 11'sd-623, 13'sd-2664}},
{{12'sd-1659, 11'sd676, 10'sd-418}, {13'sd-2310, 10'sd373, 11'sd-615}, {11'sd-760, 10'sd419, 9'sd-215}},
{{11'sd-680, 11'sd819, 12'sd1032}, {13'sd2066, 10'sd-371, 10'sd-448}, {13'sd-2135, 10'sd-379, 8'sd-70}},
{{9'sd254, 9'sd-142, 13'sd-2300}, {12'sd1277, 12'sd1044, 12'sd1051}, {12'sd1418, 8'sd-120, 10'sd-458}},
{{12'sd-1082, 10'sd-419, 13'sd-2431}, {12'sd-1583, 13'sd2245, 9'sd-207}, {13'sd2290, 11'sd-1006, 12'sd-1743}},
{{8'sd-68, 11'sd560, 13'sd-2194}, {13'sd2090, 13'sd-2659, 13'sd-2829}, {13'sd2331, 13'sd-2817, 13'sd-2796}},
{{12'sd1974, 12'sd-1343, 12'sd1345}, {13'sd-2074, 13'sd-3026, 11'sd743}, {12'sd1163, 10'sd436, 12'sd1406}},
{{12'sd-1624, 11'sd-880, 12'sd-1525}, {9'sd150, 12'sd-1427, 10'sd-385}, {11'sd791, 12'sd1201, 12'sd-1805}},
{{10'sd-349, 10'sd-290, 13'sd2236}, {11'sd619, 9'sd152, 12'sd-1325}, {12'sd-1784, 13'sd-2493, 12'sd1827}},
{{11'sd-714, 12'sd-1771, 7'sd40}, {11'sd-839, 11'sd694, 13'sd-3176}, {12'sd1526, 12'sd-1251, 11'sd-740}},
{{12'sd1185, 7'sd-51, 13'sd2289}, {8'sd-97, 8'sd101, 12'sd-1039}, {11'sd-805, 13'sd-2135, 13'sd-2481}},
{{10'sd358, 5'sd15, 12'sd-1889}, {11'sd-731, 12'sd1049, 9'sd-143}, {13'sd2512, 12'sd1345, 12'sd-1925}},
{{12'sd1269, 10'sd-493, 11'sd831}, {4'sd-6, 9'sd190, 11'sd-744}, {10'sd327, 11'sd-549, 12'sd1223}},
{{13'sd3028, 12'sd-1291, 11'sd-516}, {13'sd2675, 13'sd2262, 10'sd-402}, {11'sd-656, 10'sd-264, 10'sd-277}},
{{11'sd842, 5'sd-14, 12'sd-1432}, {10'sd282, 12'sd-1236, 13'sd3253}, {13'sd2855, 10'sd-441, 12'sd1840}},
{{13'sd-2768, 10'sd258, 12'sd-1302}, {13'sd-2142, 12'sd-1946, 13'sd-2077}, {12'sd1521, 12'sd-1599, 12'sd-1560}},
{{13'sd-2631, 13'sd-2192, 12'sd-1329}, {12'sd-1824, 12'sd1310, 13'sd2910}, {13'sd3506, 12'sd1473, 14'sd7080}},
{{13'sd2526, 12'sd-1206, 13'sd2067}, {9'sd-170, 9'sd129, 12'sd-1554}, {12'sd1570, 12'sd-1118, 10'sd302}},
{{12'sd1231, 11'sd-547, 10'sd-354}, {11'sd-899, 13'sd-2123, 13'sd-2417}, {13'sd3093, 11'sd1004, 10'sd489}},
{{11'sd-649, 11'sd-663, 9'sd-138}, {10'sd-415, 13'sd2435, 13'sd-2094}, {11'sd-884, 10'sd393, 11'sd669}},
{{13'sd3030, 8'sd116, 12'sd1536}, {12'sd-1994, 12'sd1221, 12'sd-1436}, {13'sd-2270, 13'sd-2725, 13'sd-2276}},
{{12'sd-1333, 11'sd-998, 12'sd-1781}, {13'sd-2918, 12'sd1311, 11'sd-678}, {13'sd-2078, 12'sd1503, 11'sd-557}},
{{12'sd1232, 12'sd1537, 11'sd-664}, {9'sd129, 12'sd-1702, 9'sd201}, {10'sd453, 10'sd-492, 11'sd532}},
{{11'sd808, 12'sd1345, 12'sd1358}, {13'sd2467, 12'sd-1629, 7'sd45}, {11'sd881, 11'sd819, 12'sd-1240}},
{{13'sd-2494, 12'sd-1172, 12'sd1685}, {13'sd2087, 12'sd1937, 12'sd-1396}, {12'sd1228, 11'sd836, 10'sd-479}},
{{13'sd2300, 12'sd-1617, 12'sd-1314}, {12'sd1652, 12'sd-1566, 13'sd2284}, {10'sd-385, 13'sd-4032, 12'sd1300}},
{{13'sd2264, 12'sd1930, 13'sd2278}, {10'sd488, 11'sd950, 13'sd2213}, {12'sd-1276, 12'sd-1940, 12'sd-1195}},
{{12'sd-1091, 11'sd567, 12'sd1445}, {10'sd257, 10'sd484, 13'sd3405}, {13'sd-3816, 9'sd-141, 12'sd1119}},
{{11'sd957, 11'sd-914, 13'sd-2672}, {10'sd-261, 10'sd-353, 12'sd-1073}, {12'sd1160, 12'sd-2018, 9'sd236}},
{{13'sd2828, 11'sd848, 13'sd3662}, {11'sd-808, 11'sd666, 13'sd2855}, {12'sd-1928, 10'sd-430, 9'sd180}},
{{12'sd1704, 12'sd1853, 12'sd1768}, {10'sd-333, 11'sd-671, 12'sd1150}, {11'sd602, 10'sd-309, 8'sd-111}},
{{13'sd-2919, 12'sd-1665, 11'sd758}, {10'sd366, 10'sd262, 10'sd441}, {11'sd977, 10'sd-371, 13'sd2633}},
{{12'sd1489, 12'sd1772, 13'sd-2350}, {10'sd-500, 8'sd71, 10'sd-315}, {12'sd1740, 9'sd172, 12'sd-1561}},
{{11'sd1021, 12'sd1580, 12'sd-1146}, {12'sd1389, 13'sd-2414, 13'sd2067}, {12'sd1123, 10'sd-398, 12'sd-1416}},
{{13'sd2183, 13'sd2488, 13'sd-2440}, {11'sd731, 12'sd-1127, 12'sd-1244}, {12'sd1426, 10'sd-396, 12'sd1024}},
{{11'sd606, 11'sd996, 11'sd667}, {12'sd-2018, 11'sd696, 13'sd-2138}, {11'sd-741, 12'sd-1799, 12'sd-1869}},
{{11'sd-883, 7'sd-38, 10'sd-306}, {12'sd1317, 12'sd1239, 10'sd321}, {12'sd-1088, 12'sd-1105, 12'sd-1621}}},
{
{{12'sd-1445, 12'sd-1300, 13'sd-2219}, {13'sd2315, 10'sd307, 7'sd52}, {12'sd1515, 11'sd949, 12'sd-1766}},
{{12'sd-1561, 10'sd-464, 12'sd-2046}, {13'sd-2378, 13'sd-2520, 12'sd-1738}, {11'sd-963, 12'sd-1221, 8'sd102}},
{{11'sd875, 10'sd293, 11'sd789}, {12'sd1940, 13'sd2239, 12'sd-1897}, {12'sd1355, 11'sd-790, 11'sd-764}},
{{13'sd2273, 10'sd-344, 13'sd2572}, {13'sd2526, 10'sd-409, 9'sd244}, {13'sd-2053, 12'sd1314, 9'sd-192}},
{{13'sd2140, 7'sd41, 11'sd-611}, {11'sd928, 7'sd-40, 11'sd-572}, {11'sd-764, 13'sd-2357, 10'sd309}},
{{12'sd1080, 11'sd801, 13'sd2174}, {13'sd-2416, 11'sd811, 12'sd1268}, {11'sd-649, 13'sd2921, 10'sd-286}},
{{11'sd-734, 12'sd-1740, 11'sd987}, {12'sd1599, 10'sd395, 11'sd1000}, {13'sd2506, 12'sd-1167, 10'sd-440}},
{{12'sd1113, 13'sd2876, 10'sd392}, {12'sd-1940, 13'sd2402, 10'sd454}, {8'sd70, 10'sd-281, 12'sd-1758}},
{{13'sd2322, 13'sd-2535, 13'sd2261}, {10'sd264, 12'sd-1569, 12'sd1718}, {10'sd-485, 12'sd1880, 10'sd317}},
{{12'sd1229, 12'sd1182, 12'sd2042}, {13'sd2665, 12'sd-1793, 11'sd553}, {7'sd-53, 10'sd423, 13'sd2415}},
{{12'sd1933, 12'sd-1889, 8'sd-74}, {13'sd-2400, 13'sd-2112, 11'sd-638}, {12'sd-1838, 12'sd-1542, 12'sd-1028}},
{{13'sd2728, 12'sd-1790, 10'sd430}, {12'sd1610, 13'sd2437, 10'sd-335}, {12'sd-1078, 11'sd676, 12'sd1727}},
{{8'sd-112, 12'sd1097, 12'sd-1293}, {13'sd-2833, 12'sd-1973, 11'sd537}, {12'sd-1791, 10'sd-414, 12'sd-1521}},
{{10'sd-425, 12'sd1961, 11'sd-733}, {12'sd1414, 12'sd-1301, 12'sd1024}, {9'sd-152, 11'sd-982, 13'sd-2773}},
{{10'sd368, 9'sd-128, 12'sd-1710}, {12'sd1697, 13'sd3954, 13'sd2479}, {13'sd3492, 13'sd3010, 11'sd669}},
{{12'sd1769, 11'sd850, 12'sd2034}, {10'sd400, 12'sd-1677, 9'sd-174}, {13'sd-2335, 12'sd1109, 11'sd924}},
{{10'sd-398, 10'sd-276, 10'sd306}, {12'sd1680, 11'sd543, 12'sd1188}, {9'sd-200, 13'sd-2742, 13'sd-2867}},
{{11'sd822, 13'sd-2825, 13'sd-2309}, {13'sd-2543, 10'sd349, 12'sd-1733}, {12'sd1608, 12'sd-1977, 12'sd-1331}},
{{5'sd13, 13'sd2198, 13'sd2367}, {12'sd1278, 11'sd-660, 13'sd-2283}, {13'sd-2131, 12'sd-1730, 12'sd1585}},
{{10'sd475, 12'sd1491, 13'sd-2150}, {12'sd-1961, 10'sd-401, 12'sd-1696}, {13'sd2291, 12'sd-1055, 13'sd-2712}},
{{12'sd1789, 12'sd1482, 11'sd-1005}, {13'sd-2124, 12'sd-1814, 10'sd397}, {9'sd-196, 12'sd1708, 10'sd481}},
{{10'sd430, 13'sd2436, 12'sd-1508}, {10'sd309, 13'sd2104, 12'sd-1066}, {12'sd-1260, 11'sd-1004, 11'sd-858}},
{{10'sd-313, 13'sd-2849, 12'sd-2006}, {12'sd-1159, 13'sd-2329, 13'sd2446}, {11'sd573, 12'sd-1977, 13'sd-2159}},
{{12'sd1619, 12'sd1932, 12'sd-1711}, {12'sd-1716, 13'sd2176, 12'sd1668}, {12'sd-1990, 1'sd0, 5'sd-10}},
{{10'sd484, 10'sd470, 12'sd-1757}, {12'sd1207, 12'sd-2005, 12'sd1452}, {12'sd1522, 13'sd-2154, 10'sd-257}},
{{13'sd2175, 10'sd341, 12'sd-1623}, {12'sd-1502, 11'sd889, 10'sd391}, {13'sd-2212, 12'sd-1422, 10'sd384}},
{{12'sd2022, 2'sd1, 13'sd2617}, {13'sd2124, 13'sd2222, 11'sd-878}, {8'sd-76, 13'sd-2486, 13'sd-2315}},
{{11'sd917, 13'sd-2648, 11'sd-1004}, {13'sd2976, 12'sd-1275, 12'sd1672}, {13'sd2809, 10'sd-421, 13'sd2351}},
{{13'sd2188, 12'sd-1238, 13'sd2799}, {13'sd3001, 13'sd-2316, 11'sd524}, {12'sd1264, 11'sd704, 12'sd-1393}},
{{11'sd-602, 12'sd1609, 12'sd-1991}, {13'sd2162, 11'sd604, 13'sd-2148}, {13'sd-2169, 12'sd-1475, 12'sd1133}},
{{13'sd-2488, 10'sd392, 11'sd-538}, {13'sd2688, 8'sd111, 13'sd-2201}, {10'sd339, 13'sd-2525, 12'sd1730}},
{{11'sd-845, 12'sd-1711, 10'sd268}, {12'sd-1371, 12'sd1109, 13'sd2881}, {13'sd-2527, 10'sd258, 10'sd-397}},
{{11'sd-1016, 11'sd909, 12'sd1047}, {13'sd-2403, 10'sd480, 12'sd-1224}, {12'sd1938, 13'sd2447, 11'sd913}},
{{12'sd2038, 13'sd2570, 13'sd2563}, {12'sd1784, 10'sd-465, 12'sd1124}, {12'sd1190, 13'sd2288, 11'sd948}},
{{11'sd871, 12'sd-1628, 12'sd-1302}, {10'sd470, 12'sd-1554, 13'sd-2131}, {12'sd-2011, 10'sd415, 13'sd-2385}},
{{11'sd-1000, 12'sd1823, 13'sd-2303}, {12'sd1492, 11'sd-545, 9'sd-233}, {10'sd483, 11'sd586, 12'sd-1869}},
{{12'sd1808, 12'sd-2011, 12'sd1170}, {11'sd-983, 13'sd3381, 12'sd-1257}, {11'sd-835, 12'sd1892, 11'sd-753}},
{{10'sd403, 11'sd-782, 13'sd-2509}, {13'sd-2055, 12'sd1562, 13'sd-2250}, {12'sd-1633, 10'sd-319, 13'sd-2718}},
{{11'sd872, 12'sd2044, 12'sd1380}, {12'sd-1249, 11'sd-700, 11'sd-887}, {11'sd-777, 11'sd528, 12'sd1749}},
{{12'sd1906, 12'sd1640, 12'sd-2047}, {11'sd-790, 11'sd-730, 10'sd405}, {8'sd120, 11'sd945, 13'sd2550}},
{{13'sd-2185, 11'sd782, 13'sd-2661}, {12'sd-1577, 11'sd-757, 8'sd99}, {13'sd-2258, 11'sd955, 13'sd-2084}},
{{13'sd-2934, 12'sd1308, 12'sd1661}, {11'sd-796, 12'sd-1471, 11'sd-893}, {11'sd-998, 13'sd2116, 12'sd1957}},
{{12'sd2012, 13'sd2735, 12'sd-1332}, {8'sd-100, 13'sd3006, 12'sd1691}, {11'sd-582, 13'sd2855, 12'sd-1267}},
{{12'sd-1567, 8'sd99, 12'sd-1851}, {13'sd-2535, 12'sd1270, 13'sd-3348}, {13'sd-2345, 12'sd-1415, 13'sd-3465}},
{{12'sd-1883, 12'sd-1223, 12'sd1619}, {11'sd-515, 12'sd1117, 11'sd-689}, {13'sd-2576, 10'sd-277, 11'sd739}},
{{12'sd-1731, 13'sd-2329, 12'sd1223}, {10'sd261, 12'sd-1842, 12'sd1645}, {12'sd-1254, 8'sd-88, 12'sd1942}},
{{11'sd-725, 12'sd1539, 13'sd2591}, {12'sd1036, 11'sd789, 12'sd2044}, {13'sd-2978, 12'sd-1699, 9'sd-178}},
{{12'sd-1467, 12'sd-1248, 9'sd142}, {13'sd-2299, 13'sd2214, 12'sd1964}, {12'sd1166, 7'sd-56, 11'sd680}},
{{12'sd1687, 11'sd-622, 12'sd1280}, {12'sd1274, 13'sd2756, 12'sd-1252}, {13'sd-2322, 11'sd-989, 13'sd2276}},
{{13'sd2397, 12'sd1290, 10'sd-367}, {12'sd-1307, 12'sd-1240, 13'sd2844}, {12'sd1044, 13'sd2210, 11'sd-641}},
{{12'sd1860, 12'sd-1203, 11'sd514}, {13'sd2431, 8'sd-102, 3'sd-3}, {10'sd431, 11'sd982, 11'sd683}},
{{12'sd1889, 11'sd513, 12'sd-1159}, {11'sd-836, 10'sd-264, 13'sd-2475}, {12'sd-1907, 12'sd-1755, 13'sd2248}},
{{11'sd609, 12'sd1595, 12'sd-1337}, {12'sd2047, 12'sd1542, 9'sd133}, {11'sd755, 11'sd-726, 9'sd241}},
{{13'sd-2365, 12'sd1187, 13'sd-2606}, {12'sd1670, 11'sd-766, 10'sd323}, {12'sd2014, 13'sd2165, 10'sd346}},
{{13'sd2308, 11'sd795, 12'sd1275}, {13'sd2691, 10'sd-319, 13'sd-2389}, {11'sd532, 13'sd2247, 12'sd1613}},
{{13'sd2401, 10'sd-275, 10'sd-300}, {12'sd-1942, 12'sd-1941, 12'sd-1202}, {11'sd925, 12'sd1683, 9'sd183}},
{{13'sd-2122, 9'sd-142, 11'sd-532}, {10'sd332, 11'sd-566, 12'sd-1741}, {12'sd1655, 12'sd1088, 13'sd2583}},
{{11'sd932, 12'sd-1865, 13'sd-2111}, {13'sd2206, 12'sd1200, 10'sd349}, {10'sd300, 13'sd-2053, 12'sd-1171}},
{{12'sd1674, 9'sd-157, 13'sd-2247}, {9'sd-199, 13'sd-2413, 12'sd-1631}, {11'sd-845, 11'sd715, 13'sd-2076}},
{{13'sd2185, 7'sd35, 13'sd2487}, {12'sd-1988, 13'sd-2294, 11'sd854}, {9'sd-135, 12'sd1807, 12'sd1771}},
{{11'sd857, 12'sd1113, 12'sd1294}, {12'sd1417, 10'sd507, 13'sd-2757}, {11'sd-717, 10'sd-382, 10'sd258}},
{{12'sd1145, 13'sd2361, 13'sd-2506}, {10'sd-410, 11'sd972, 11'sd-619}, {12'sd1271, 10'sd499, 9'sd-168}},
{{11'sd989, 11'sd-781, 12'sd-1488}, {12'sd1682, 12'sd1434, 12'sd-1281}, {13'sd2500, 13'sd-2099, 13'sd2321}},
{{12'sd-1297, 11'sd523, 12'sd1290}, {12'sd-1825, 13'sd3670, 11'sd888}, {12'sd-1427, 11'sd-766, 12'sd-1149}}},
{
{{13'sd-2841, 11'sd-792, 12'sd-1921}, {11'sd-943, 11'sd529, 10'sd299}, {10'sd-350, 12'sd-1230, 10'sd-261}},
{{13'sd3358, 12'sd1779, 12'sd1211}, {9'sd-225, 12'sd-1781, 13'sd-2124}, {10'sd-270, 12'sd2001, 13'sd-2511}},
{{13'sd3106, 12'sd1776, 13'sd2630}, {13'sd-2497, 11'sd-534, 12'sd-1320}, {11'sd-903, 13'sd-2215, 9'sd-238}},
{{11'sd-733, 13'sd-2965, 11'sd692}, {13'sd2129, 12'sd-1604, 13'sd2106}, {11'sd695, 9'sd-145, 11'sd922}},
{{13'sd3400, 8'sd120, 12'sd-1408}, {12'sd1170, 11'sd883, 11'sd840}, {12'sd1492, 11'sd555, 13'sd-2173}},
{{12'sd-2017, 14'sd-4385, 14'sd-4839}, {11'sd762, 11'sd762, 10'sd297}, {12'sd1560, 8'sd-122, 11'sd545}},
{{11'sd626, 11'sd-747, 14'sd-5026}, {11'sd606, 10'sd460, 12'sd-1330}, {13'sd-2081, 12'sd-1997, 14'sd-5293}},
{{11'sd-946, 12'sd-1195, 12'sd1205}, {10'sd-438, 12'sd1878, 12'sd-1251}, {12'sd-1787, 11'sd574, 12'sd-1850}},
{{10'sd-314, 11'sd-1001, 12'sd-1680}, {9'sd-129, 9'sd251, 12'sd1152}, {13'sd-2820, 11'sd-540, 10'sd256}},
{{11'sd-599, 12'sd1487, 13'sd-2512}, {12'sd-1971, 11'sd-773, 12'sd-1643}, {13'sd-2807, 11'sd949, 10'sd425}},
{{13'sd3860, 11'sd-773, 12'sd-1092}, {11'sd-804, 12'sd-1986, 9'sd148}, {13'sd-3038, 11'sd742, 13'sd-2113}},
{{10'sd334, 11'sd514, 12'sd1231}, {13'sd3024, 10'sd-261, 13'sd-2328}, {9'sd192, 12'sd1106, 11'sd-898}},
{{12'sd1835, 12'sd1607, 12'sd-1836}, {13'sd2472, 12'sd1570, 13'sd-2477}, {11'sd1008, 9'sd-206, 13'sd-3001}},
{{13'sd2569, 12'sd1828, 12'sd2004}, {11'sd699, 11'sd934, 12'sd1726}, {11'sd-720, 10'sd-384, 12'sd1782}},
{{12'sd1526, 12'sd1226, 13'sd-2208}, {13'sd-2341, 12'sd1174, 14'sd-4177}, {6'sd-25, 14'sd4103, 11'sd-992}},
{{5'sd-9, 13'sd2633, 11'sd935}, {12'sd1334, 13'sd2297, 13'sd3330}, {10'sd462, 12'sd-1827, 13'sd-2426}},
{{13'sd-3279, 10'sd-369, 13'sd-2482}, {13'sd2056, 11'sd-1008, 12'sd1077}, {12'sd1964, 13'sd2872, 12'sd-1397}},
{{13'sd3523, 12'sd1316, 11'sd992}, {13'sd3114, 13'sd2294, 11'sd769}, {13'sd2319, 11'sd658, 11'sd638}},
{{10'sd-347, 13'sd2227, 12'sd1648}, {12'sd1544, 12'sd1730, 10'sd-476}, {12'sd-1186, 13'sd2354, 12'sd-1213}},
{{8'sd118, 13'sd-2364, 13'sd-2226}, {12'sd-1905, 13'sd-2124, 10'sd-316}, {12'sd1404, 13'sd2067, 13'sd2304}},
{{13'sd-2334, 11'sd584, 12'sd1944}, {13'sd-3065, 11'sd730, 13'sd-2338}, {12'sd-1678, 11'sd-636, 11'sd-976}},
{{13'sd-3187, 13'sd-2184, 13'sd-2124}, {9'sd176, 10'sd364, 11'sd-521}, {13'sd2643, 11'sd-697, 13'sd3146}},
{{12'sd1120, 12'sd-1535, 11'sd946}, {12'sd1863, 12'sd1623, 13'sd2739}, {13'sd-2057, 12'sd1640, 13'sd-2302}},
{{13'sd-2892, 13'sd-2586, 12'sd-1806}, {11'sd-638, 11'sd585, 11'sd927}, {12'sd-1067, 13'sd2536, 13'sd3113}},
{{12'sd1159, 12'sd-1568, 11'sd920}, {13'sd2282, 13'sd-2505, 7'sd-40}, {13'sd2677, 12'sd-1124, 12'sd-1093}},
{{12'sd-1073, 10'sd-335, 13'sd2105}, {10'sd-380, 12'sd1107, 12'sd1344}, {12'sd-1360, 9'sd-201, 13'sd-3584}},
{{11'sd580, 10'sd418, 9'sd151}, {12'sd-1077, 11'sd-826, 11'sd-933}, {10'sd282, 12'sd-1418, 13'sd-4081}},
{{13'sd3033, 12'sd1366, 10'sd432}, {13'sd2554, 12'sd-1176, 8'sd85}, {13'sd-2250, 13'sd-2049, 13'sd-2953}},
{{11'sd649, 12'sd1347, 12'sd1961}, {11'sd-561, 13'sd2570, 10'sd-353}, {13'sd-2333, 12'sd2002, 12'sd1923}},
{{13'sd2260, 12'sd-1560, 12'sd1233}, {13'sd2096, 12'sd1719, 10'sd462}, {12'sd-1931, 12'sd-1146, 13'sd2827}},
{{13'sd-2163, 12'sd1482, 12'sd-1553}, {11'sd810, 13'sd-2240, 11'sd-523}, {12'sd-1226, 12'sd1615, 13'sd-2161}},
{{9'sd-233, 11'sd-864, 13'sd-2751}, {12'sd1874, 11'sd-937, 12'sd-1529}, {10'sd-381, 10'sd511, 9'sd160}},
{{13'sd-2955, 13'sd-2199, 11'sd-913}, {8'sd-97, 11'sd-947, 11'sd-751}, {12'sd1290, 13'sd-2550, 12'sd1474}},
{{13'sd2882, 11'sd521, 11'sd707}, {13'sd2366, 10'sd385, 11'sd940}, {13'sd2360, 11'sd954, 13'sd3527}},
{{12'sd1930, 11'sd870, 11'sd920}, {12'sd1944, 11'sd-869, 11'sd732}, {12'sd-1472, 12'sd1439, 12'sd1360}},
{{13'sd-2375, 13'sd-2276, 12'sd-1280}, {10'sd-501, 12'sd-1214, 12'sd-1996}, {12'sd-1791, 12'sd1860, 11'sd655}},
{{12'sd-1067, 11'sd-953, 12'sd-1115}, {12'sd-2001, 8'sd-122, 12'sd1504}, {12'sd1867, 11'sd550, 14'sd4757}},
{{11'sd-601, 13'sd2594, 11'sd817}, {12'sd-1995, 12'sd-1632, 12'sd-1434}, {13'sd-2592, 11'sd861, 11'sd861}},
{{7'sd-52, 11'sd-695, 10'sd390}, {12'sd-1347, 12'sd1386, 11'sd-575}, {10'sd501, 12'sd-1225, 12'sd1769}},
{{8'sd79, 13'sd-2080, 12'sd-1062}, {11'sd728, 12'sd-1213, 13'sd-2406}, {13'sd-2260, 12'sd1456, 11'sd744}},
{{13'sd-2080, 12'sd1672, 12'sd-1729}, {8'sd73, 13'sd2485, 12'sd-1349}, {12'sd1044, 10'sd302, 12'sd1476}},
{{13'sd4043, 12'sd1342, 13'sd2703}, {12'sd-1842, 12'sd-1169, 12'sd1575}, {14'sd-4628, 14'sd-5940, 13'sd-2628}},
{{7'sd49, 12'sd1820, 12'sd1101}, {13'sd2202, 8'sd-110, 11'sd817}, {13'sd-2166, 10'sd466, 12'sd-1116}},
{{14'sd5425, 13'sd2253, 13'sd3537}, {14'sd4598, 13'sd-2062, 11'sd-1004}, {13'sd3002, 13'sd-3327, 13'sd-3545}},
{{11'sd944, 9'sd175, 12'sd-1658}, {11'sd-879, 13'sd2145, 13'sd-2513}, {12'sd-1079, 10'sd473, 11'sd-1000}},
{{12'sd-1621, 10'sd296, 13'sd-3004}, {12'sd-1998, 13'sd-2986, 11'sd954}, {13'sd2744, 12'sd1558, 12'sd1993}},
{{11'sd-966, 9'sd-234, 13'sd-2123}, {11'sd-557, 12'sd1054, 7'sd51}, {5'sd-12, 10'sd420, 12'sd-1214}},
{{13'sd3219, 11'sd-795, 11'sd-823}, {12'sd-1867, 11'sd-1014, 11'sd-586}, {13'sd3293, 12'sd1564, 12'sd1225}},
{{13'sd2592, 12'sd1884, 7'sd-46}, {8'sd121, 12'sd1694, 12'sd-1796}, {12'sd1623, 13'sd2377, 12'sd1359}},
{{14'sd-5945, 13'sd-3439, 12'sd-1286}, {11'sd-611, 13'sd-3108, 13'sd2829}, {12'sd-1747, 13'sd4031, 10'sd503}},
{{11'sd-941, 12'sd1970, 9'sd210}, {12'sd1999, 11'sd-775, 12'sd1797}, {12'sd-1214, 11'sd696, 12'sd1801}},
{{10'sd-294, 9'sd136, 12'sd-1818}, {12'sd-1360, 12'sd-1084, 13'sd-2162}, {13'sd-2255, 12'sd1523, 6'sd-19}},
{{12'sd1381, 12'sd-1876, 13'sd-2089}, {10'sd281, 12'sd-1963, 9'sd214}, {9'sd169, 13'sd-2350, 11'sd-948}},
{{11'sd646, 13'sd-2171, 9'sd-161}, {12'sd2043, 12'sd-1221, 11'sd-972}, {12'sd-1704, 12'sd1924, 13'sd-2282}},
{{12'sd-1908, 13'sd-2537, 13'sd-3244}, {13'sd2341, 12'sd-2023, 13'sd-2281}, {14'sd-5131, 12'sd-1893, 14'sd-5744}},
{{13'sd-3653, 12'sd-1770, 12'sd-1784}, {7'sd-56, 12'sd-1229, 12'sd-1671}, {12'sd-1489, 13'sd-2100, 13'sd3180}},
{{11'sd739, 12'sd-1510, 10'sd310}, {13'sd-2649, 12'sd-1510, 10'sd426}, {13'sd-3389, 13'sd-2084, 14'sd-5693}},
{{13'sd2681, 13'sd2359, 10'sd-286}, {13'sd2178, 12'sd-1752, 12'sd1388}, {11'sd-532, 12'sd-1218, 12'sd1883}},
{{13'sd2833, 11'sd561, 12'sd-1619}, {11'sd566, 13'sd2704, 12'sd1070}, {13'sd-3237, 13'sd-3057, 9'sd-252}},
{{12'sd1462, 12'sd-1446, 8'sd85}, {12'sd1810, 14'sd4139, 11'sd-884}, {12'sd-1335, 11'sd-527, 12'sd-2045}},
{{10'sd-342, 13'sd-2127, 11'sd612}, {12'sd1564, 12'sd-1758, 12'sd1134}, {10'sd491, 12'sd1720, 13'sd3370}},
{{9'sd-231, 13'sd-2129, 10'sd-288}, {12'sd1877, 10'sd286, 12'sd-1715}, {12'sd-1955, 12'sd-1061, 12'sd-1439}},
{{11'sd-952, 13'sd-2488, 13'sd2076}, {13'sd2255, 12'sd-1513, 13'sd2153}, {12'sd-1921, 9'sd-220, 12'sd1029}},
{{9'sd-148, 13'sd-3395, 6'sd-21}, {11'sd864, 12'sd1308, 12'sd-1314}, {12'sd1758, 13'sd3224, 11'sd-934}}},
{
{{13'sd-3061, 13'sd-2421, 12'sd1513}, {11'sd-641, 11'sd-735, 12'sd1822}, {11'sd872, 10'sd440, 12'sd1896}},
{{13'sd2777, 7'sd60, 11'sd515}, {11'sd-963, 12'sd1238, 11'sd-699}, {12'sd1428, 11'sd512, 12'sd1455}},
{{12'sd1772, 12'sd-1676, 12'sd-1092}, {9'sd-156, 13'sd-2564, 10'sd329}, {11'sd-598, 11'sd-563, 12'sd-1590}},
{{13'sd-2517, 12'sd-1708, 12'sd-1549}, {9'sd-217, 9'sd146, 13'sd2615}, {12'sd1631, 10'sd-420, 13'sd-2116}},
{{13'sd2619, 13'sd2191, 13'sd2679}, {13'sd3842, 12'sd-1945, 12'sd1190}, {13'sd-3259, 13'sd-2628, 9'sd183}},
{{13'sd3001, 12'sd1736, 11'sd994}, {13'sd2862, 12'sd-1622, 13'sd2853}, {10'sd-317, 13'sd-2079, 13'sd2241}},
{{13'sd2197, 13'sd-3429, 13'sd3302}, {12'sd1502, 13'sd-2712, 12'sd-1653}, {13'sd4076, 12'sd1350, 13'sd2958}},
{{12'sd-1463, 13'sd-2401, 12'sd1284}, {12'sd1279, 13'sd2138, 13'sd2992}, {11'sd670, 11'sd-527, 12'sd1870}},
{{10'sd307, 12'sd1962, 9'sd-136}, {13'sd2189, 12'sd-1448, 13'sd-2809}, {12'sd1304, 12'sd1337, 11'sd-692}},
{{7'sd59, 12'sd1098, 13'sd2434}, {11'sd-961, 13'sd2875, 12'sd-1865}, {12'sd1653, 12'sd1661, 10'sd401}},
{{13'sd-2702, 11'sd-697, 12'sd-1156}, {13'sd-2784, 9'sd253, 12'sd1344}, {13'sd-3386, 9'sd156, 12'sd-1463}},
{{13'sd2295, 8'sd82, 13'sd2778}, {10'sd358, 13'sd2107, 10'sd-389}, {13'sd-2597, 9'sd-206, 13'sd-3053}},
{{12'sd-1656, 10'sd-314, 11'sd660}, {12'sd-1629, 11'sd1021, 12'sd1224}, {12'sd-1476, 12'sd1089, 13'sd-2166}},
{{12'sd1290, 12'sd1321, 9'sd-255}, {11'sd-689, 11'sd-738, 13'sd2638}, {10'sd456, 13'sd-2856, 13'sd-2519}},
{{12'sd-1089, 13'sd-2285, 10'sd323}, {11'sd581, 11'sd668, 12'sd1578}, {12'sd-1923, 11'sd-794, 12'sd-1162}},
{{12'sd1498, 13'sd2426, 12'sd1970}, {11'sd-602, 12'sd-1424, 13'sd-3039}, {12'sd1376, 10'sd291, 12'sd-1270}},
{{10'sd-448, 10'sd-502, 12'sd-1531}, {12'sd1896, 12'sd1834, 12'sd-1551}, {12'sd-1492, 9'sd-246, 11'sd674}},
{{11'sd830, 11'sd654, 13'sd2343}, {12'sd1303, 12'sd-1591, 12'sd1131}, {13'sd-2389, 11'sd-1003, 12'sd1374}},
{{12'sd1953, 13'sd2864, 12'sd-1425}, {12'sd1921, 12'sd-1106, 13'sd2369}, {11'sd990, 10'sd462, 12'sd-1819}},
{{11'sd954, 12'sd-1853, 11'sd653}, {13'sd2903, 10'sd-325, 11'sd-922}, {13'sd2742, 12'sd-1142, 11'sd-772}},
{{12'sd-1214, 8'sd67, 12'sd-1358}, {12'sd-2036, 13'sd-2775, 11'sd548}, {11'sd-892, 11'sd-1022, 12'sd2019}},
{{10'sd-264, 12'sd-1075, 12'sd1395}, {11'sd872, 12'sd1348, 12'sd-1607}, {11'sd719, 13'sd-2140, 11'sd860}},
{{13'sd3649, 12'sd-1069, 12'sd1639}, {13'sd2696, 1'sd0, 11'sd794}, {12'sd1596, 13'sd-2382, 12'sd1645}},
{{12'sd-1751, 12'sd-1875, 12'sd-1071}, {11'sd-969, 12'sd1105, 11'sd-642}, {11'sd-819, 11'sd740, 11'sd1004}},
{{11'sd655, 13'sd2472, 3'sd3}, {10'sd-283, 12'sd-1123, 12'sd1447}, {11'sd-979, 12'sd-1344, 13'sd-2455}},
{{13'sd-2638, 10'sd403, 12'sd-1718}, {12'sd-1406, 11'sd741, 13'sd2583}, {10'sd-424, 13'sd-2635, 12'sd1428}},
{{13'sd-2863, 13'sd-2238, 13'sd-2890}, {13'sd-4013, 12'sd1284, 12'sd1847}, {12'sd-1810, 10'sd310, 13'sd2557}},
{{13'sd-2096, 12'sd-1354, 13'sd2540}, {13'sd-2696, 8'sd79, 12'sd1088}, {12'sd-1748, 12'sd1718, 12'sd2023}},
{{7'sd-36, 12'sd1581, 10'sd272}, {12'sd1386, 12'sd-1140, 13'sd-2643}, {10'sd469, 12'sd-1413, 12'sd-1737}},
{{12'sd-1727, 13'sd2380, 12'sd-1387}, {12'sd1548, 11'sd634, 12'sd-1234}, {10'sd-470, 11'sd-959, 13'sd3058}},
{{10'sd-493, 11'sd-565, 11'sd876}, {10'sd-451, 13'sd2230, 12'sd1879}, {13'sd2333, 10'sd-488, 12'sd1353}},
{{9'sd136, 12'sd-1906, 12'sd-1303}, {13'sd-2432, 13'sd-2686, 10'sd-434}, {13'sd2721, 12'sd1146, 11'sd1005}},
{{12'sd-1903, 10'sd-495, 12'sd-1998}, {9'sd185, 10'sd331, 13'sd-2475}, {11'sd873, 10'sd-385, 12'sd-1484}},
{{11'sd-1009, 13'sd2507, 13'sd-2184}, {12'sd1642, 12'sd-1248, 13'sd-3040}, {12'sd1278, 11'sd515, 12'sd1940}},
{{7'sd45, 11'sd-944, 10'sd325}, {12'sd-1377, 6'sd-31, 10'sd293}, {13'sd-2578, 12'sd1704, 10'sd338}},
{{13'sd3330, 12'sd-2006, 10'sd272}, {11'sd909, 12'sd-1042, 12'sd-1664}, {7'sd32, 11'sd516, 12'sd-1962}},
{{14'sd-4576, 14'sd-4298, 12'sd-1451}, {12'sd1666, 10'sd282, 13'sd-2097}, {13'sd3366, 11'sd735, 11'sd-588}},
{{11'sd-684, 9'sd-152, 12'sd-1466}, {13'sd3353, 13'sd2637, 8'sd104}, {11'sd654, 12'sd1734, 12'sd1249}},
{{11'sd617, 11'sd-675, 12'sd1070}, {10'sd-434, 11'sd695, 12'sd-1470}, {8'sd78, 12'sd-1809, 13'sd-2389}},
{{10'sd396, 13'sd-2113, 12'sd2002}, {12'sd1555, 12'sd1298, 12'sd1471}, {11'sd-741, 10'sd500, 12'sd2047}},
{{14'sd4496, 12'sd1027, 11'sd590}, {13'sd2109, 11'sd849, 8'sd104}, {9'sd-191, 12'sd1965, 10'sd353}},
{{12'sd-1579, 13'sd-2460, 10'sd486}, {12'sd1991, 12'sd1231, 13'sd-2300}, {13'sd-2092, 13'sd-2685, 11'sd538}},
{{12'sd-1518, 12'sd1279, 10'sd-290}, {9'sd233, 12'sd1451, 11'sd570}, {12'sd-1124, 12'sd1312, 11'sd-616}},
{{13'sd-2184, 13'sd-2885, 9'sd213}, {11'sd802, 12'sd-1841, 13'sd-2314}, {13'sd-2893, 11'sd-749, 14'sd-5051}},
{{13'sd-2303, 9'sd-156, 12'sd-1950}, {12'sd-1860, 9'sd-222, 13'sd2486}, {12'sd-1861, 12'sd-1024, 12'sd-1566}},
{{10'sd450, 13'sd-2480, 13'sd2382}, {12'sd1281, 12'sd1519, 11'sd561}, {10'sd458, 10'sd-304, 12'sd1512}},
{{12'sd-1554, 13'sd-2382, 8'sd78}, {11'sd692, 13'sd-2227, 11'sd-806}, {11'sd-642, 12'sd1114, 12'sd1344}},
{{12'sd-1531, 9'sd-244, 12'sd-1845}, {13'sd-2261, 12'sd-1984, 12'sd1102}, {5'sd11, 12'sd-2039, 12'sd1026}},
{{11'sd-858, 11'sd-705, 13'sd2755}, {13'sd-2516, 10'sd350, 12'sd1640}, {12'sd1984, 12'sd1512, 13'sd2937}},
{{3'sd2, 11'sd-1017, 13'sd-3391}, {12'sd1135, 10'sd447, 12'sd1528}, {13'sd-2167, 10'sd457, 12'sd1369}},
{{10'sd443, 12'sd1209, 12'sd1376}, {12'sd-1757, 12'sd1453, 11'sd-939}, {13'sd2216, 12'sd1929, 12'sd-1150}},
{{12'sd-1618, 12'sd-1131, 13'sd-2785}, {11'sd542, 9'sd211, 10'sd364}, {9'sd-188, 11'sd675, 13'sd2643}},
{{12'sd1617, 10'sd436, 12'sd-1168}, {4'sd7, 13'sd2115, 12'sd1687}, {13'sd-3295, 13'sd-2672, 12'sd-1271}},
{{11'sd-1009, 12'sd1156, 11'sd-900}, {12'sd-1035, 13'sd-2412, 13'sd-2420}, {12'sd-1337, 12'sd1639, 13'sd-2278}},
{{13'sd-2672, 12'sd-1228, 10'sd-395}, {11'sd929, 10'sd-490, 13'sd2208}, {12'sd1806, 13'sd3195, 13'sd2119}},
{{13'sd-2152, 13'sd-2706, 13'sd-2543}, {12'sd-1525, 11'sd635, 13'sd-2067}, {12'sd-1144, 12'sd-1128, 12'sd1782}},
{{12'sd-1070, 12'sd1966, 13'sd-2278}, {12'sd1502, 12'sd-2032, 10'sd-301}, {13'sd-3032, 13'sd-4025, 14'sd-4204}},
{{10'sd-289, 12'sd1968, 13'sd2493}, {13'sd3036, 11'sd618, 13'sd-2657}, {12'sd1190, 11'sd-683, 13'sd-3090}},
{{7'sd55, 12'sd1940, 10'sd358}, {11'sd588, 12'sd-1599, 13'sd2296}, {5'sd9, 12'sd-1818, 12'sd1962}},
{{12'sd1777, 13'sd3917, 13'sd2276}, {12'sd1101, 13'sd-2084, 12'sd1334}, {13'sd2632, 12'sd1143, 13'sd2660}},
{{12'sd1090, 12'sd1217, 13'sd-2401}, {12'sd1751, 11'sd705, 12'sd1507}, {12'sd-1243, 12'sd1719, 13'sd-2118}},
{{10'sd499, 13'sd2557, 13'sd-2273}, {12'sd1312, 12'sd-2045, 13'sd2768}, {12'sd-1096, 12'sd1762, 11'sd889}},
{{11'sd914, 12'sd1255, 12'sd-1732}, {12'sd1286, 12'sd-1049, 10'sd300}, {13'sd-2571, 13'sd2342, 12'sd-1784}},
{{12'sd-1353, 13'sd-2907, 11'sd870}, {13'sd-2856, 13'sd-2334, 12'sd-1281}, {7'sd-48, 11'sd1023, 13'sd2453}}},
{
{{11'sd-797, 13'sd-2099, 11'sd852}, {11'sd-862, 12'sd1407, 11'sd990}, {11'sd-605, 11'sd681, 12'sd1230}},
{{12'sd1501, 13'sd-3121, 12'sd-1609}, {13'sd-2542, 10'sd-475, 11'sd-636}, {13'sd-2064, 11'sd772, 12'sd-1900}},
{{12'sd-1135, 9'sd141, 12'sd-1621}, {12'sd2030, 10'sd-488, 13'sd2238}, {12'sd-1482, 12'sd-1957, 12'sd-1696}},
{{11'sd-732, 12'sd-1543, 13'sd2559}, {12'sd1495, 12'sd-1698, 12'sd1318}, {13'sd2702, 12'sd-1725, 12'sd-1875}},
{{13'sd-2433, 12'sd1962, 13'sd2345}, {13'sd-3471, 10'sd-400, 13'sd-2174}, {14'sd-4096, 12'sd-1420, 13'sd-4002}},
{{9'sd166, 13'sd2186, 13'sd3026}, {13'sd-2419, 13'sd-2682, 12'sd1168}, {13'sd-2072, 13'sd-2298, 12'sd1205}},
{{10'sd330, 12'sd1509, 13'sd3420}, {11'sd820, 10'sd377, 13'sd2890}, {13'sd2454, 11'sd-593, 9'sd-218}},
{{11'sd744, 12'sd1799, 9'sd240}, {13'sd-2274, 11'sd-717, 11'sd-789}, {13'sd-2234, 6'sd-25, 11'sd808}},
{{13'sd2481, 13'sd-2108, 11'sd987}, {12'sd1434, 12'sd1416, 13'sd-2748}, {12'sd-1520, 13'sd2313, 10'sd334}},
{{12'sd1936, 12'sd-1683, 12'sd-2012}, {12'sd1429, 12'sd-1934, 12'sd-1445}, {13'sd3497, 13'sd2906, 11'sd571}},
{{6'sd27, 12'sd-1926, 10'sd-354}, {12'sd-1645, 12'sd1257, 12'sd-1421}, {13'sd2546, 12'sd1640, 9'sd-182}},
{{12'sd-1709, 13'sd2482, 9'sd187}, {10'sd444, 12'sd-1289, 10'sd-312}, {13'sd-2401, 13'sd2205, 13'sd-2239}},
{{11'sd-869, 12'sd-1950, 13'sd-3301}, {11'sd906, 12'sd-1957, 11'sd1018}, {12'sd1636, 13'sd2319, 13'sd-2053}},
{{11'sd883, 9'sd222, 10'sd-441}, {10'sd329, 12'sd-1615, 13'sd-2570}, {12'sd1301, 12'sd1616, 13'sd-2393}},
{{12'sd-1432, 9'sd196, 11'sd641}, {12'sd1507, 13'sd3037, 13'sd3582}, {13'sd3334, 6'sd30, 10'sd-300}},
{{12'sd-1735, 9'sd251, 12'sd-1749}, {12'sd-1136, 12'sd-1676, 12'sd1071}, {11'sd-618, 13'sd-2603, 11'sd-865}},
{{12'sd1865, 13'sd2501, 10'sd440}, {9'sd-186, 13'sd2411, 13'sd2390}, {12'sd-1945, 12'sd-1332, 13'sd-2815}},
{{12'sd-1151, 8'sd-74, 12'sd-1816}, {13'sd2256, 12'sd-1491, 10'sd383}, {13'sd2128, 12'sd1612, 10'sd509}},
{{12'sd-1634, 11'sd630, 12'sd-1781}, {11'sd1019, 12'sd-1424, 9'sd-189}, {12'sd-1387, 13'sd2053, 8'sd-79}},
{{13'sd-2578, 13'sd-2242, 12'sd1369}, {9'sd161, 13'sd2353, 12'sd-1408}, {10'sd-283, 12'sd-2022, 12'sd1207}},
{{12'sd-1081, 12'sd1897, 13'sd2819}, {12'sd-1113, 13'sd2148, 11'sd-896}, {12'sd1487, 11'sd906, 11'sd868}},
{{11'sd-1006, 13'sd-2375, 12'sd1368}, {11'sd706, 9'sd179, 11'sd-875}, {13'sd-2285, 8'sd90, 7'sd59}},
{{13'sd2603, 10'sd-453, 13'sd-2591}, {13'sd-2321, 12'sd1190, 12'sd-1095}, {12'sd1682, 12'sd1049, 10'sd-295}},
{{10'sd-407, 13'sd-2131, 13'sd-2069}, {10'sd347, 10'sd-445, 12'sd1061}, {11'sd1006, 11'sd935, 12'sd-1126}},
{{13'sd-2402, 10'sd-294, 11'sd-599}, {10'sd421, 10'sd-354, 7'sd42}, {13'sd-2622, 13'sd-2985, 12'sd-1579}},
{{11'sd-703, 11'sd-947, 11'sd-850}, {12'sd-1736, 12'sd-1281, 11'sd591}, {9'sd224, 13'sd-2512, 12'sd1089}},
{{12'sd-1902, 12'sd-1639, 13'sd-2165}, {13'sd-3719, 13'sd-2275, 13'sd-2517}, {10'sd265, 12'sd1060, 4'sd-4}},
{{12'sd-1151, 12'sd-1581, 12'sd1083}, {11'sd-773, 11'sd891, 10'sd478}, {13'sd-2324, 9'sd-186, 12'sd1746}},
{{10'sd-424, 12'sd1351, 12'sd1895}, {12'sd1553, 9'sd131, 13'sd3231}, {12'sd-1997, 12'sd1591, 10'sd-351}},
{{13'sd-2917, 11'sd-1000, 12'sd1309}, {11'sd816, 11'sd-664, 13'sd-2468}, {12'sd-1251, 12'sd1981, 13'sd-2162}},
{{10'sd-402, 12'sd-1188, 12'sd1910}, {13'sd2528, 12'sd-1520, 12'sd1469}, {12'sd-1924, 13'sd-2299, 12'sd-1207}},
{{12'sd-1135, 9'sd195, 13'sd2270}, {13'sd2359, 10'sd441, 11'sd974}, {12'sd1636, 11'sd-769, 13'sd3317}},
{{12'sd1878, 12'sd-1275, 13'sd2238}, {12'sd-1454, 13'sd-2691, 12'sd1793}, {12'sd-1747, 10'sd-463, 12'sd-1671}},
{{10'sd326, 13'sd-2562, 11'sd928}, {12'sd-1753, 13'sd-2172, 12'sd-1920}, {12'sd-1165, 12'sd2016, 12'sd-1872}},
{{10'sd-368, 12'sd1943, 12'sd1546}, {13'sd-2228, 11'sd645, 11'sd950}, {12'sd-1062, 12'sd-1025, 13'sd-2307}},
{{9'sd152, 11'sd869, 13'sd2905}, {11'sd-618, 12'sd1027, 10'sd-370}, {12'sd1805, 12'sd1812, 9'sd146}},
{{13'sd-3820, 13'sd2199, 13'sd2666}, {10'sd-421, 13'sd2491, 12'sd1909}, {9'sd-178, 13'sd-2079, 12'sd1165}},
{{12'sd-1751, 12'sd-1511, 12'sd1564}, {12'sd2031, 12'sd-1917, 13'sd-2731}, {10'sd362, 11'sd913, 11'sd655}},
{{13'sd-2054, 11'sd922, 12'sd-2037}, {13'sd-2259, 13'sd2307, 12'sd1952}, {12'sd1226, 11'sd534, 4'sd7}},
{{11'sd832, 12'sd1037, 11'sd1002}, {13'sd-2141, 11'sd-513, 12'sd1950}, {12'sd1110, 10'sd-499, 9'sd-143}},
{{12'sd-1528, 13'sd2437, 11'sd695}, {9'sd-165, 11'sd629, 11'sd851}, {13'sd-2386, 10'sd288, 10'sd405}},
{{11'sd830, 11'sd611, 12'sd1375}, {11'sd648, 10'sd-363, 13'sd-2450}, {13'sd2985, 12'sd1867, 10'sd-406}},
{{10'sd-388, 12'sd-1469, 12'sd1230}, {8'sd114, 12'sd1936, 11'sd930}, {13'sd2410, 13'sd2492, 11'sd-783}},
{{7'sd-61, 11'sd-645, 13'sd-3185}, {12'sd-1829, 13'sd2209, 10'sd430}, {14'sd-5719, 14'sd-4119, 10'sd-267}},
{{13'sd-2709, 12'sd-1495, 13'sd2454}, {13'sd2081, 11'sd668, 12'sd1236}, {12'sd1476, 11'sd1016, 12'sd1834}},
{{13'sd2522, 13'sd2505, 13'sd2760}, {12'sd-1528, 11'sd669, 12'sd1816}, {13'sd-3310, 11'sd823, 11'sd-815}},
{{14'sd-4291, 10'sd281, 11'sd-625}, {8'sd-120, 8'sd-79, 13'sd2342}, {11'sd1001, 12'sd1334, 13'sd3144}},
{{11'sd-711, 12'sd-1875, 13'sd3322}, {13'sd-2825, 12'sd-1634, 12'sd-2031}, {10'sd476, 13'sd2309, 10'sd290}},
{{10'sd-495, 8'sd118, 12'sd1773}, {12'sd-1466, 13'sd2751, 12'sd-1404}, {12'sd-1109, 12'sd-1538, 13'sd2349}},
{{13'sd-2620, 12'sd-1482, 12'sd-1772}, {12'sd-1239, 11'sd-701, 13'sd3449}, {10'sd387, 12'sd1517, 11'sd-711}},
{{13'sd-2079, 12'sd-1367, 11'sd519}, {12'sd1671, 12'sd1838, 12'sd1039}, {12'sd-1686, 13'sd-2680, 10'sd-357}},
{{8'sd78, 11'sd1021, 13'sd2580}, {12'sd1444, 11'sd-681, 12'sd1280}, {12'sd1173, 13'sd2231, 13'sd-2210}},
{{13'sd2921, 12'sd1224, 12'sd-1978}, {11'sd-667, 12'sd1741, 13'sd2650}, {10'sd410, 11'sd581, 12'sd1126}},
{{11'sd-941, 10'sd-285, 12'sd-1121}, {11'sd815, 13'sd-2308, 8'sd87}, {12'sd-1225, 12'sd1523, 13'sd2515}},
{{13'sd-2139, 13'sd-2811, 13'sd-2462}, {13'sd-2261, 13'sd-2283, 13'sd-3850}, {12'sd-1622, 13'sd2096, 13'sd2592}},
{{9'sd185, 12'sd1500, 9'sd-211}, {9'sd219, 13'sd2693, 13'sd2478}, {13'sd-2451, 11'sd996, 12'sd-1677}},
{{12'sd1048, 11'sd647, 10'sd275}, {12'sd1315, 13'sd-2276, 12'sd-1098}, {11'sd538, 11'sd-954, 13'sd-2670}},
{{10'sd269, 8'sd119, 12'sd-1716}, {9'sd189, 13'sd-2927, 13'sd-2997}, {11'sd-940, 11'sd-610, 12'sd1204}},
{{12'sd-1673, 12'sd1481, 13'sd-2120}, {12'sd1736, 10'sd414, 12'sd1300}, {13'sd2506, 13'sd2519, 12'sd1218}},
{{9'sd226, 13'sd3105, 13'sd3863}, {13'sd-2768, 12'sd-1547, 13'sd-2070}, {13'sd-2243, 8'sd85, 13'sd2723}},
{{13'sd-2824, 12'sd1635, 11'sd-1020}, {12'sd1258, 13'sd-2242, 12'sd1566}, {12'sd-1608, 12'sd-1855, 12'sd1192}},
{{12'sd1175, 12'sd-1686, 13'sd2420}, {11'sd-758, 11'sd-536, 13'sd-2365}, {12'sd1221, 12'sd-1341, 12'sd-1751}},
{{11'sd586, 13'sd-2977, 13'sd-2932}, {11'sd-833, 12'sd1075, 10'sd269}, {11'sd953, 11'sd-769, 10'sd396}},
{{13'sd3599, 11'sd-512, 13'sd4034}, {13'sd3141, 13'sd2894, 13'sd2520}, {13'sd2270, 12'sd1993, 13'sd2597}}},
{
{{12'sd1113, 12'sd1782, 13'sd2174}, {13'sd-2770, 10'sd-337, 13'sd-2063}, {12'sd-1944, 12'sd-1614, 8'sd-73}},
{{11'sd-802, 11'sd987, 10'sd277}, {10'sd-419, 12'sd-1679, 12'sd-1936}, {7'sd35, 12'sd-1391, 13'sd-2434}},
{{12'sd-1877, 12'sd1933, 13'sd2065}, {12'sd-1695, 12'sd-1907, 11'sd802}, {13'sd2084, 11'sd-678, 10'sd-468}},
{{13'sd-2090, 9'sd235, 11'sd587}, {12'sd-1531, 12'sd1067, 10'sd402}, {13'sd-2454, 10'sd267, 12'sd1492}},
{{14'sd-4135, 13'sd-2112, 11'sd880}, {13'sd-2303, 13'sd2270, 9'sd150}, {3'sd-3, 9'sd-182, 11'sd-901}},
{{12'sd-1633, 13'sd-3992, 13'sd-2834}, {13'sd-3693, 12'sd1106, 9'sd-163}, {13'sd2328, 13'sd-2939, 12'sd-1744}},
{{13'sd-3324, 9'sd167, 13'sd-4036}, {11'sd948, 12'sd1774, 11'sd681}, {13'sd-3169, 12'sd-1294, 13'sd-3518}},
{{12'sd1121, 12'sd-1445, 12'sd1077}, {13'sd-2049, 10'sd-407, 11'sd-801}, {10'sd285, 12'sd1471, 10'sd308}},
{{13'sd-2709, 12'sd-1147, 10'sd-278}, {13'sd-3030, 13'sd2369, 10'sd-445}, {11'sd980, 9'sd-195, 12'sd-1881}},
{{6'sd-20, 11'sd879, 12'sd-1557}, {12'sd-1289, 10'sd338, 10'sd315}, {12'sd2043, 12'sd1737, 13'sd-2930}},
{{12'sd1592, 13'sd2928, 9'sd-213}, {11'sd-947, 12'sd1863, 12'sd-1930}, {11'sd734, 13'sd-2302, 8'sd-73}},
{{10'sd417, 12'sd-1947, 9'sd-189}, {13'sd-2057, 12'sd-1853, 12'sd1642}, {13'sd-2679, 12'sd-1911, 13'sd2766}},
{{12'sd1839, 12'sd-1378, 11'sd742}, {12'sd1456, 13'sd2664, 9'sd132}, {11'sd955, 8'sd106, 12'sd1623}},
{{6'sd-26, 9'sd213, 12'sd-1681}, {10'sd324, 10'sd-339, 9'sd-158}, {11'sd-882, 12'sd-1766, 12'sd1735}},
{{13'sd-3991, 12'sd1899, 13'sd4021}, {7'sd-39, 13'sd3706, 13'sd3936}, {12'sd-1145, 11'sd1010, 14'sd4848}},
{{12'sd1978, 13'sd2294, 12'sd-1121}, {12'sd1145, 11'sd-872, 11'sd-885}, {12'sd-1411, 10'sd375, 10'sd-399}},
{{6'sd-26, 13'sd2379, 10'sd-431}, {10'sd378, 11'sd-612, 12'sd1591}, {10'sd325, 11'sd-914, 10'sd-267}},
{{12'sd-1460, 13'sd-2131, 10'sd302}, {9'sd222, 13'sd-2551, 12'sd-1383}, {12'sd-1485, 13'sd2251, 13'sd2235}},
{{13'sd2332, 12'sd-1217, 11'sd846}, {12'sd1317, 13'sd2507, 13'sd-2963}, {11'sd735, 12'sd-1332, 13'sd-2146}},
{{8'sd82, 13'sd-2366, 13'sd-2146}, {11'sd965, 13'sd-2581, 10'sd413}, {12'sd1155, 13'sd-2426, 12'sd-1890}},
{{11'sd-1013, 11'sd-570, 12'sd1209}, {12'sd-1976, 9'sd-131, 12'sd-1814}, {11'sd-788, 11'sd991, 12'sd1432}},
{{10'sd-386, 9'sd-200, 12'sd1360}, {10'sd-377, 13'sd-2430, 13'sd-2538}, {13'sd2262, 13'sd-2092, 8'sd-98}},
{{13'sd-2626, 12'sd1122, 11'sd-938}, {13'sd2345, 12'sd-1514, 12'sd-1750}, {13'sd2874, 12'sd1419, 12'sd-1579}},
{{12'sd1784, 9'sd-200, 12'sd1778}, {13'sd-2231, 11'sd-852, 10'sd486}, {10'sd-269, 12'sd-1972, 10'sd-506}},
{{13'sd2614, 13'sd-2291, 13'sd-2655}, {13'sd-2195, 10'sd461, 12'sd1785}, {12'sd1707, 6'sd30, 12'sd1324}},
{{12'sd1126, 11'sd-513, 12'sd1657}, {12'sd1445, 13'sd2845, 7'sd52}, {11'sd608, 12'sd-1149, 12'sd-1780}},
{{14'sd6374, 12'sd1658, 12'sd-1368}, {11'sd753, 11'sd719, 12'sd-1507}, {11'sd569, 14'sd-5065, 13'sd-3529}},
{{11'sd851, 11'sd879, 12'sd-1091}, {11'sd-699, 8'sd117, 12'sd1315}, {10'sd-476, 13'sd-2317, 10'sd341}},
{{12'sd1802, 13'sd2798, 11'sd519}, {11'sd-534, 11'sd819, 13'sd3835}, {12'sd1875, 10'sd-471, 13'sd2746}},
{{12'sd1974, 13'sd-2553, 10'sd349}, {13'sd2607, 12'sd-1758, 13'sd-2244}, {9'sd201, 13'sd-2087, 11'sd-911}},
{{12'sd-1388, 11'sd599, 11'sd-567}, {8'sd-98, 9'sd-145, 13'sd-2964}, {11'sd520, 13'sd2442, 12'sd1275}},
{{12'sd-1567, 12'sd-1609, 13'sd2069}, {12'sd1196, 12'sd1224, 12'sd2022}, {11'sd532, 12'sd1597, 8'sd91}},
{{13'sd-2676, 12'sd-1933, 10'sd319}, {12'sd-1623, 12'sd-1597, 12'sd1944}, {13'sd2116, 13'sd-2223, 12'sd1438}},
{{13'sd-3034, 10'sd-352, 11'sd-653}, {12'sd-1457, 12'sd1344, 12'sd1387}, {12'sd-1222, 12'sd-1038, 12'sd-1704}},
{{12'sd-1789, 12'sd1483, 13'sd-2283}, {12'sd1225, 8'sd-101, 9'sd228}, {12'sd1764, 12'sd1128, 13'sd-2078}},
{{12'sd1993, 13'sd-2995, 12'sd2002}, {13'sd-2165, 11'sd806, 12'sd-1593}, {12'sd-1935, 12'sd-1583, 13'sd2606}},
{{13'sd3554, 11'sd537, 13'sd3568}, {12'sd1623, 9'sd-193, 12'sd1316}, {11'sd-754, 12'sd-1175, 12'sd1906}},
{{13'sd2317, 12'sd1538, 11'sd-930}, {11'sd-776, 12'sd-1768, 13'sd-3192}, {13'sd2433, 5'sd12, 9'sd217}},
{{12'sd-1773, 11'sd-878, 13'sd-2637}, {10'sd502, 12'sd-1746, 12'sd-1727}, {11'sd-648, 13'sd-2213, 12'sd-2024}},
{{12'sd-1137, 12'sd1662, 11'sd-846}, {12'sd-1092, 9'sd-134, 12'sd-1640}, {10'sd-371, 12'sd-1461, 8'sd-100}},
{{12'sd1125, 13'sd-2327, 13'sd-3583}, {13'sd2121, 13'sd-2779, 12'sd-1043}, {12'sd-1931, 13'sd-3045, 12'sd-2017}},
{{12'sd-1276, 12'sd-1086, 12'sd1263}, {13'sd3386, 12'sd1334, 13'sd2717}, {12'sd1029, 11'sd807, 13'sd2134}},
{{11'sd700, 11'sd638, 11'sd-625}, {12'sd1610, 13'sd2209, 11'sd977}, {12'sd1551, 12'sd-2014, 12'sd1793}},
{{14'sd8092, 14'sd6122, 12'sd1295}, {14'sd7311, 11'sd913, 14'sd-4758}, {13'sd2938, 12'sd1735, 13'sd-2905}},
{{10'sd-477, 12'sd1441, 12'sd2016}, {11'sd-861, 13'sd2579, 13'sd2162}, {12'sd-1529, 10'sd320, 8'sd96}},
{{12'sd1063, 12'sd1889, 11'sd698}, {12'sd1945, 13'sd2778, 10'sd507}, {12'sd1247, 12'sd-1784, 10'sd439}},
{{12'sd1747, 13'sd3063, 13'sd2446}, {13'sd2953, 11'sd659, 12'sd-1791}, {12'sd-1520, 12'sd1065, 13'sd-2230}},
{{11'sd-682, 12'sd1440, 12'sd-1968}, {13'sd2325, 10'sd-359, 12'sd1584}, {12'sd1679, 12'sd1994, 11'sd892}},
{{11'sd-719, 11'sd603, 12'sd-1033}, {13'sd-3558, 9'sd-202, 12'sd-1161}, {13'sd-3412, 12'sd-1405, 12'sd-1317}},
{{12'sd-1319, 13'sd-2092, 11'sd-751}, {12'sd1877, 13'sd-2914, 6'sd-21}, {12'sd1589, 12'sd1964, 13'sd2272}},
{{12'sd-1977, 11'sd-562, 11'sd991}, {11'sd-784, 12'sd2029, 11'sd851}, {12'sd1250, 13'sd-2296, 13'sd3112}},
{{10'sd-301, 12'sd-2010, 13'sd-2646}, {12'sd-1098, 12'sd-1672, 13'sd2203}, {12'sd-1593, 12'sd-1889, 9'sd230}},
{{12'sd2031, 6'sd-21, 12'sd-1078}, {12'sd-2041, 13'sd2732, 12'sd-1638}, {11'sd514, 11'sd-628, 11'sd-628}},
{{12'sd1942, 13'sd-2081, 12'sd-1350}, {12'sd-1938, 11'sd-640, 12'sd1670}, {8'sd75, 11'sd-572, 12'sd-1137}},
{{13'sd-2319, 13'sd-2138, 10'sd-269}, {13'sd2879, 12'sd2019, 13'sd-2928}, {10'sd-458, 12'sd1223, 11'sd715}},
{{13'sd-2716, 10'sd488, 11'sd-649}, {13'sd-2385, 12'sd1399, 11'sd-892}, {11'sd669, 10'sd-309, 13'sd2278}},
{{14'sd4157, 13'sd-2692, 13'sd2517}, {13'sd2089, 9'sd204, 9'sd-176}, {13'sd3139, 13'sd2491, 11'sd694}},
{{12'sd-1887, 13'sd2997, 13'sd2426}, {12'sd-2001, 10'sd-304, 12'sd-1126}, {9'sd-198, 12'sd-1797, 13'sd-2250}},
{{11'sd-637, 11'sd639, 13'sd-2594}, {12'sd-1082, 10'sd301, 9'sd236}, {12'sd-1470, 12'sd1997, 11'sd-850}},
{{13'sd-3519, 10'sd-507, 10'sd-386}, {12'sd-1499, 11'sd611, 13'sd2939}, {13'sd-2470, 11'sd790, 10'sd-274}},
{{12'sd1378, 13'sd-3116, 13'sd2353}, {11'sd856, 13'sd-2589, 11'sd856}, {13'sd2580, 12'sd1109, 13'sd2051}},
{{13'sd-2147, 13'sd2210, 11'sd672}, {11'sd-728, 10'sd397, 12'sd1851}, {12'sd-1478, 12'sd-1635, 12'sd1894}},
{{13'sd3315, 12'sd1234, 13'sd2403}, {11'sd-779, 11'sd1023, 13'sd-3180}, {13'sd2365, 11'sd725, 13'sd-2304}},
{{12'sd1743, 12'sd-1463, 10'sd-469}, {8'sd-114, 12'sd-1677, 10'sd334}, {12'sd-1392, 13'sd2533, 12'sd-1897}}},
{
{{12'sd-1876, 8'sd-91, 13'sd-2266}, {6'sd-29, 13'sd-2096, 12'sd-1235}, {11'sd988, 12'sd-1100, 12'sd-1708}},
{{12'sd1437, 12'sd1976, 12'sd1605}, {11'sd-521, 11'sd-932, 12'sd-1521}, {10'sd413, 11'sd886, 11'sd524}},
{{12'sd-1324, 9'sd137, 10'sd-453}, {13'sd-2815, 12'sd-1995, 12'sd1054}, {8'sd83, 10'sd471, 12'sd1791}},
{{13'sd-2402, 13'sd2353, 13'sd-2526}, {10'sd417, 11'sd1021, 13'sd-2243}, {12'sd-1732, 10'sd499, 12'sd1271}},
{{10'sd361, 10'sd-438, 14'sd-6006}, {13'sd-2562, 10'sd-301, 13'sd-2949}, {13'sd-3177, 12'sd1805, 13'sd-2236}},
{{13'sd3556, 11'sd696, 13'sd3983}, {13'sd-2073, 13'sd3520, 12'sd1115}, {12'sd-1565, 13'sd2953, 11'sd806}},
{{11'sd-940, 12'sd1381, 12'sd-1183}, {11'sd-973, 12'sd1730, 13'sd-2175}, {13'sd-2595, 14'sd5451, 12'sd1361}},
{{11'sd577, 13'sd2655, 12'sd1962}, {12'sd-1762, 11'sd926, 12'sd-1329}, {12'sd1969, 9'sd240, 12'sd1537}},
{{12'sd-1587, 12'sd1241, 12'sd1345}, {12'sd-2031, 11'sd-994, 13'sd-2196}, {11'sd610, 13'sd-2419, 12'sd1567}},
{{11'sd805, 11'sd649, 11'sd-814}, {13'sd-3565, 13'sd-2325, 13'sd-2386}, {11'sd692, 13'sd2105, 12'sd-1283}},
{{13'sd-2084, 10'sd-297, 11'sd660}, {13'sd2368, 8'sd89, 13'sd2818}, {13'sd-2177, 13'sd-2103, 12'sd-1964}},
{{13'sd3188, 12'sd1089, 12'sd1098}, {12'sd-1830, 13'sd-2306, 13'sd-2930}, {9'sd203, 11'sd638, 12'sd1242}},
{{14'sd-4256, 12'sd-1678, 12'sd1148}, {11'sd-1010, 11'sd922, 12'sd-1315}, {7'sd60, 11'sd546, 12'sd-1316}},
{{11'sd549, 10'sd-470, 12'sd-1440}, {11'sd581, 12'sd-1397, 11'sd582}, {12'sd-1033, 13'sd2137, 11'sd526}},
{{13'sd3963, 10'sd-425, 15'sd-8999}, {12'sd1143, 14'sd-4356, 13'sd-3980}, {12'sd-2019, 13'sd2224, 11'sd526}},
{{10'sd282, 12'sd1625, 7'sd55}, {12'sd-1431, 12'sd-1580, 13'sd-3017}, {12'sd1806, 11'sd786, 12'sd1897}},
{{11'sd-930, 13'sd-3118, 9'sd181}, {12'sd1281, 13'sd2436, 12'sd1627}, {12'sd-1343, 7'sd-38, 12'sd1064}},
{{9'sd191, 8'sd78, 12'sd1061}, {11'sd973, 12'sd1726, 12'sd1673}, {13'sd-3054, 11'sd737, 7'sd-46}},
{{13'sd-2823, 9'sd174, 11'sd-784}, {12'sd1545, 12'sd-1028, 12'sd1172}, {12'sd-1358, 13'sd2316, 11'sd-677}},
{{11'sd1010, 12'sd-2004, 9'sd167}, {13'sd2912, 11'sd620, 12'sd-1192}, {10'sd-330, 10'sd-354, 11'sd819}},
{{8'sd-85, 12'sd1839, 13'sd-2512}, {10'sd333, 12'sd1680, 9'sd-145}, {11'sd884, 8'sd-124, 12'sd-1061}},
{{11'sd612, 10'sd-511, 8'sd-113}, {12'sd1085, 8'sd90, 12'sd-1919}, {12'sd-1657, 11'sd892, 7'sd-43}},
{{10'sd-487, 11'sd-526, 12'sd-1568}, {12'sd-1319, 10'sd-444, 13'sd-2774}, {13'sd-3062, 10'sd481, 12'sd-1419}},
{{13'sd-2260, 10'sd-491, 12'sd1074}, {9'sd-129, 13'sd-2167, 12'sd1982}, {13'sd-2136, 12'sd1946, 12'sd1753}},
{{13'sd-2180, 13'sd-2860, 10'sd-270}, {12'sd-1323, 11'sd844, 8'sd71}, {9'sd169, 12'sd1941, 9'sd133}},
{{7'sd-56, 13'sd2514, 12'sd1228}, {11'sd-903, 12'sd-1738, 8'sd-70}, {13'sd-2213, 13'sd-2208, 13'sd-2861}},
{{11'sd647, 14'sd5185, 14'sd8018}, {12'sd1944, 12'sd1634, 14'sd5154}, {13'sd3271, 9'sd-232, 9'sd186}},
{{12'sd1719, 13'sd2643, 13'sd-3912}, {13'sd-2160, 12'sd1551, 13'sd-2959}, {10'sd-475, 10'sd353, 12'sd1430}},
{{12'sd1495, 6'sd-25, 11'sd929}, {11'sd763, 12'sd1073, 12'sd-1221}, {12'sd1824, 10'sd-367, 8'sd-88}},
{{11'sd959, 11'sd-556, 14'sd4498}, {13'sd2826, 13'sd2742, 13'sd3743}, {13'sd2742, 12'sd1205, 11'sd-637}},
{{12'sd-1056, 12'sd-1114, 10'sd-388}, {12'sd1900, 12'sd-1363, 13'sd2256}, {12'sd-1220, 12'sd1300, 13'sd2418}},
{{13'sd-2539, 12'sd-1775, 13'sd-2175}, {10'sd-347, 12'sd1396, 10'sd-282}, {13'sd2173, 11'sd-955, 13'sd-2351}},
{{12'sd1139, 13'sd-2990, 10'sd-415}, {11'sd849, 12'sd-1220, 12'sd-1340}, {12'sd2018, 10'sd-391, 12'sd-1344}},
{{11'sd-897, 12'sd1397, 13'sd2476}, {13'sd-2189, 12'sd-1784, 13'sd-2466}, {13'sd-2459, 12'sd1553, 13'sd2678}},
{{14'sd5438, 13'sd2241, 12'sd-1053}, {14'sd4414, 11'sd-711, 13'sd2201}, {12'sd1216, 12'sd1464, 10'sd-273}},
{{12'sd1169, 13'sd-2581, 11'sd827}, {10'sd-491, 13'sd-3342, 10'sd394}, {12'sd1702, 12'sd1246, 12'sd-1480}},
{{14'sd4174, 13'sd3218, 13'sd2309}, {14'sd6748, 12'sd1321, 13'sd2474}, {14'sd7775, 14'sd4598, 12'sd1370}},
{{10'sd464, 13'sd2614, 13'sd-2512}, {13'sd2373, 12'sd1286, 12'sd1943}, {13'sd-2559, 13'sd2628, 11'sd-909}},
{{12'sd-1938, 11'sd987, 12'sd1535}, {11'sd-760, 12'sd-1714, 12'sd1484}, {12'sd1744, 9'sd-177, 13'sd-2958}},
{{12'sd1200, 13'sd-2911, 8'sd-121}, {13'sd2295, 12'sd-1844, 12'sd-1285}, {10'sd-314, 13'sd-2352, 12'sd-1237}},
{{13'sd4037, 12'sd1421, 12'sd1959}, {13'sd3155, 13'sd3070, 12'sd1056}, {11'sd759, 11'sd526, 12'sd1440}},
{{13'sd-2810, 13'sd-2820, 10'sd-443}, {12'sd-1714, 9'sd237, 12'sd1626}, {13'sd-2174, 9'sd235, 13'sd-3621}},
{{12'sd1439, 13'sd2499, 14'sd4412}, {13'sd-3539, 13'sd3450, 12'sd1884}, {11'sd-840, 13'sd2192, 12'sd1909}},
{{13'sd-3967, 10'sd-331, 12'sd-1712}, {14'sd4329, 14'sd5879, 13'sd3242}, {8'sd-109, 9'sd-241, 13'sd-2694}},
{{9'sd-163, 8'sd-81, 12'sd1889}, {12'sd-1988, 12'sd1028, 13'sd-2984}, {11'sd692, 10'sd473, 13'sd2517}},
{{12'sd2011, 12'sd-1264, 12'sd-1582}, {11'sd-532, 10'sd453, 11'sd-854}, {13'sd-2743, 9'sd131, 12'sd-1557}},
{{6'sd26, 12'sd1849, 12'sd-1943}, {13'sd2327, 10'sd476, 13'sd-2191}, {14'sd4377, 12'sd2028, 12'sd-1975}},
{{11'sd-609, 12'sd1683, 10'sd-271}, {9'sd-218, 13'sd2170, 12'sd1632}, {13'sd-2308, 9'sd-245, 12'sd-1666}},
{{13'sd3094, 11'sd969, 13'sd2377}, {10'sd320, 11'sd531, 12'sd-1711}, {14'sd4200, 11'sd810, 11'sd-1002}},
{{13'sd-2577, 13'sd-3141, 9'sd-135}, {13'sd-2198, 13'sd-2250, 13'sd-2181}, {12'sd-1954, 11'sd772, 10'sd401}},
{{14'sd4223, 12'sd1793, 12'sd-1959}, {7'sd-59, 10'sd-300, 9'sd-252}, {13'sd-3267, 11'sd-735, 8'sd127}},
{{10'sd-269, 10'sd504, 13'sd2730}, {11'sd905, 13'sd-2064, 9'sd-177}, {13'sd-2155, 12'sd1362, 13'sd-2684}},
{{9'sd-225, 12'sd-1106, 13'sd-2106}, {13'sd-2814, 11'sd-895, 6'sd27}, {12'sd-1190, 12'sd1330, 12'sd1275}},
{{12'sd1657, 9'sd-202, 13'sd-2228}, {12'sd-1564, 13'sd3000, 12'sd-2037}, {12'sd1615, 13'sd2136, 13'sd-2762}},
{{13'sd-3685, 13'sd2253, 10'sd-492}, {13'sd-4013, 11'sd792, 11'sd-750}, {8'sd117, 13'sd-3080, 11'sd552}},
{{13'sd-2273, 12'sd-1370, 12'sd-1437}, {11'sd651, 13'sd2434, 9'sd-202}, {11'sd646, 13'sd2307, 13'sd-2333}},
{{14'sd-5299, 13'sd-2719, 12'sd-1124}, {13'sd-2103, 12'sd1239, 11'sd-639}, {12'sd-1191, 14'sd-4236, 13'sd2853}},
{{10'sd260, 12'sd1369, 10'sd324}, {13'sd2282, 13'sd-3083, 12'sd1286}, {12'sd-1084, 12'sd-1710, 12'sd1253}},
{{11'sd583, 12'sd1577, 13'sd2584}, {13'sd-2781, 12'sd1109, 12'sd-1616}, {11'sd605, 12'sd1697, 11'sd-553}},
{{12'sd1258, 10'sd-361, 13'sd-3546}, {10'sd508, 10'sd-511, 14'sd-5426}, {12'sd-1846, 13'sd-2274, 12'sd-1980}},
{{12'sd1825, 13'sd-2977, 9'sd-133}, {13'sd-2282, 13'sd-2654, 10'sd452}, {9'sd-212, 9'sd176, 13'sd-2051}},
{{12'sd1929, 12'sd1058, 12'sd1393}, {11'sd827, 13'sd-2113, 13'sd-3647}, {12'sd-1074, 13'sd2055, 12'sd1171}},
{{13'sd3747, 12'sd-1298, 13'sd-2269}, {13'sd3209, 12'sd1325, 11'sd684}, {13'sd2091, 12'sd-1478, 12'sd-1738}},
{{13'sd-3517, 13'sd-2742, 13'sd-2390}, {12'sd-1935, 12'sd1530, 9'sd-212}, {13'sd3071, 12'sd1593, 12'sd1546}}},
{
{{12'sd-1619, 13'sd-2180, 13'sd2246}, {13'sd-2493, 13'sd-2516, 12'sd1977}, {13'sd2349, 12'sd-1515, 10'sd-495}},
{{12'sd-1888, 11'sd1019, 13'sd2417}, {13'sd-2542, 13'sd-2177, 11'sd589}, {11'sd-725, 12'sd-1913, 12'sd1243}},
{{11'sd-977, 13'sd2423, 11'sd952}, {12'sd-1170, 11'sd-853, 10'sd344}, {8'sd-68, 9'sd-248, 10'sd-294}},
{{12'sd-1920, 13'sd2431, 12'sd1205}, {12'sd1752, 13'sd2761, 13'sd-2536}, {11'sd-802, 12'sd1030, 9'sd-139}},
{{13'sd2576, 11'sd-973, 10'sd510}, {12'sd1226, 12'sd1177, 9'sd215}, {13'sd2566, 12'sd1293, 13'sd2359}},
{{9'sd235, 12'sd-1071, 10'sd434}, {13'sd-2317, 12'sd-1871, 13'sd-3344}, {12'sd1802, 8'sd88, 12'sd1424}},
{{12'sd-1728, 12'sd-1026, 12'sd-1335}, {12'sd1705, 10'sd493, 13'sd-2364}, {8'sd78, 9'sd-250, 12'sd1700}},
{{12'sd-1182, 13'sd2471, 11'sd557}, {10'sd321, 10'sd368, 11'sd793}, {12'sd-1318, 11'sd853, 12'sd1900}},
{{13'sd2424, 13'sd-2305, 13'sd-2720}, {12'sd-1668, 10'sd341, 13'sd2185}, {12'sd-1375, 13'sd2611, 10'sd373}},
{{13'sd-2853, 9'sd249, 12'sd-1907}, {12'sd1850, 12'sd1685, 12'sd1512}, {13'sd-2951, 13'sd2075, 11'sd520}},
{{13'sd-2721, 13'sd2098, 11'sd707}, {13'sd2136, 12'sd-1543, 10'sd494}, {11'sd-774, 9'sd230, 13'sd2129}},
{{11'sd-723, 10'sd302, 12'sd1862}, {12'sd1633, 11'sd659, 12'sd-1684}, {9'sd140, 12'sd-1866, 9'sd-162}},
{{12'sd1493, 11'sd-968, 13'sd2325}, {12'sd1538, 11'sd796, 13'sd2535}, {13'sd2377, 13'sd2324, 12'sd-1509}},
{{9'sd-241, 7'sd-38, 9'sd-171}, {12'sd1174, 12'sd-1199, 12'sd-1685}, {13'sd-2159, 11'sd709, 13'sd-2802}},
{{13'sd2579, 12'sd-1960, 5'sd15}, {7'sd-53, 13'sd2223, 11'sd729}, {13'sd2829, 13'sd2099, 13'sd3532}},
{{12'sd-1515, 13'sd2433, 11'sd680}, {13'sd-2564, 12'sd-1942, 12'sd-1531}, {12'sd-1484, 10'sd499, 11'sd825}},
{{13'sd2119, 12'sd1604, 12'sd1850}, {12'sd-1161, 12'sd-1693, 11'sd582}, {11'sd-867, 12'sd-2024, 13'sd-2293}},
{{13'sd2270, 13'sd2970, 10'sd381}, {13'sd2983, 11'sd817, 13'sd-2403}, {9'sd170, 12'sd-1644, 10'sd288}},
{{12'sd1337, 11'sd775, 13'sd-2322}, {13'sd2431, 12'sd1613, 13'sd2853}, {10'sd470, 13'sd2131, 11'sd904}},
{{12'sd-1298, 10'sd-353, 11'sd816}, {13'sd2095, 12'sd-1699, 13'sd2354}, {10'sd-357, 9'sd-223, 13'sd-2693}},
{{12'sd-1366, 13'sd-2397, 13'sd-2259}, {13'sd2906, 12'sd1207, 13'sd-2254}, {12'sd1592, 11'sd-854, 13'sd-2331}},
{{13'sd-2489, 11'sd-940, 13'sd2213}, {12'sd1968, 13'sd2398, 11'sd998}, {12'sd-1864, 11'sd966, 10'sd404}},
{{13'sd2679, 11'sd-1019, 11'sd-1009}, {12'sd-1900, 12'sd1980, 11'sd-888}, {13'sd-2853, 11'sd724, 12'sd1581}},
{{4'sd-4, 11'sd-931, 12'sd-1122}, {12'sd1603, 12'sd1302, 11'sd-823}, {12'sd1925, 10'sd264, 13'sd2538}},
{{12'sd1835, 12'sd-1473, 12'sd1120}, {10'sd369, 13'sd2517, 11'sd-565}, {12'sd1531, 13'sd-2403, 10'sd424}},
{{10'sd-273, 10'sd-448, 10'sd407}, {13'sd2273, 11'sd-596, 12'sd1327}, {12'sd1297, 13'sd-2055, 13'sd2424}},
{{13'sd2485, 12'sd1190, 12'sd1557}, {11'sd-823, 11'sd-1001, 10'sd-332}, {12'sd-1735, 10'sd-339, 12'sd1456}},
{{12'sd1582, 6'sd17, 11'sd-730}, {10'sd482, 13'sd2293, 12'sd-1476}, {13'sd3314, 13'sd3056, 12'sd-1649}},
{{11'sd910, 10'sd341, 9'sd161}, {12'sd-1063, 9'sd-195, 13'sd2748}, {12'sd-1311, 8'sd82, 11'sd844}},
{{12'sd-2038, 10'sd-265, 13'sd2676}, {11'sd-675, 10'sd483, 12'sd-1102}, {12'sd2001, 13'sd-2214, 10'sd424}},
{{10'sd276, 12'sd1246, 9'sd152}, {13'sd2094, 10'sd-427, 12'sd1534}, {13'sd-2470, 11'sd-804, 11'sd-702}},
{{13'sd-2149, 12'sd1073, 11'sd-914}, {9'sd251, 10'sd-365, 10'sd-261}, {13'sd-2247, 12'sd1812, 12'sd1526}},
{{10'sd-290, 9'sd215, 13'sd2799}, {12'sd1604, 10'sd-364, 11'sd-856}, {9'sd-205, 13'sd-2904, 12'sd1534}},
{{12'sd-1310, 12'sd-1737, 12'sd-1142}, {9'sd-242, 11'sd-736, 11'sd852}, {12'sd-1089, 12'sd1041, 10'sd422}},
{{13'sd-2613, 10'sd403, 8'sd70}, {8'sd-77, 13'sd2149, 11'sd519}, {13'sd2570, 7'sd33, 6'sd23}},
{{11'sd734, 11'sd-677, 12'sd-1601}, {5'sd10, 12'sd1102, 12'sd1938}, {13'sd-2419, 12'sd-1060, 9'sd-171}},
{{10'sd-456, 11'sd976, 11'sd631}, {12'sd-1505, 11'sd-916, 12'sd1379}, {13'sd-3225, 12'sd1889, 13'sd-2735}},
{{12'sd-1037, 13'sd-2146, 11'sd722}, {11'sd-786, 13'sd2348, 12'sd-1582}, {10'sd320, 10'sd355, 13'sd-2735}},
{{12'sd-1905, 9'sd-157, 6'sd24}, {12'sd1141, 13'sd2380, 13'sd-2385}, {9'sd231, 13'sd-2648, 11'sd837}},
{{13'sd2365, 12'sd1450, 9'sd182}, {13'sd-2088, 11'sd545, 8'sd-81}, {12'sd1066, 12'sd1902, 11'sd663}},
{{10'sd-343, 12'sd1849, 13'sd2065}, {13'sd2414, 13'sd2675, 11'sd866}, {12'sd1470, 13'sd2452, 12'sd-1649}},
{{10'sd397, 12'sd1742, 11'sd-838}, {10'sd-308, 12'sd1860, 13'sd2883}, {11'sd765, 13'sd2219, 13'sd3453}},
{{9'sd130, 13'sd2591, 10'sd-312}, {10'sd-366, 12'sd-1040, 12'sd-1180}, {9'sd160, 12'sd-1197, 13'sd3268}},
{{14'sd-4982, 11'sd-588, 14'sd-4478}, {12'sd-1836, 13'sd2652, 12'sd-1634}, {13'sd2274, 10'sd-402, 13'sd2478}},
{{12'sd-1284, 12'sd1615, 9'sd-207}, {13'sd-2216, 11'sd-660, 10'sd-313}, {10'sd435, 12'sd-1488, 13'sd-2285}},
{{12'sd-1949, 13'sd-2808, 11'sd-730}, {10'sd333, 12'sd1655, 12'sd1774}, {11'sd-905, 10'sd437, 10'sd-261}},
{{12'sd-1840, 12'sd1033, 13'sd2747}, {11'sd570, 13'sd2437, 11'sd568}, {13'sd2109, 13'sd2319, 12'sd-1893}},
{{12'sd-1529, 12'sd1167, 13'sd2556}, {12'sd-1744, 13'sd2847, 13'sd2288}, {12'sd-1741, 12'sd1231, 8'sd-113}},
{{12'sd-1676, 12'sd-1783, 12'sd-1976}, {12'sd-1990, 11'sd-686, 12'sd-1656}, {13'sd2486, 7'sd48, 12'sd1299}},
{{13'sd-2759, 12'sd-1826, 10'sd320}, {11'sd-575, 13'sd-2427, 12'sd-1747}, {12'sd1828, 9'sd189, 13'sd-2656}},
{{11'sd-764, 12'sd1311, 12'sd-1676}, {12'sd1820, 12'sd1913, 13'sd2153}, {11'sd-913, 7'sd-46, 11'sd666}},
{{10'sd258, 12'sd-1652, 12'sd-1171}, {13'sd2231, 13'sd2529, 12'sd1507}, {12'sd1310, 9'sd239, 10'sd-423}},
{{13'sd-2698, 11'sd-641, 13'sd-2587}, {13'sd-2223, 12'sd1978, 11'sd-674}, {12'sd1874, 13'sd3473, 13'sd2283}},
{{10'sd292, 13'sd-2487, 12'sd1117}, {12'sd1888, 11'sd-641, 13'sd-2308}, {11'sd-526, 12'sd-1055, 5'sd12}},
{{10'sd-288, 13'sd2654, 8'sd-103}, {13'sd3130, 12'sd-1528, 10'sd-389}, {12'sd-1866, 12'sd1481, 13'sd-2448}},
{{12'sd-1255, 13'sd-2233, 12'sd1358}, {11'sd-666, 9'sd237, 11'sd-613}, {11'sd963, 12'sd-1938, 12'sd-1231}},
{{13'sd-2137, 12'sd1183, 13'sd3036}, {14'sd4643, 11'sd850, 13'sd2071}, {14'sd5793, 13'sd3103, 13'sd3686}},
{{9'sd-148, 12'sd1248, 12'sd-1852}, {13'sd2654, 12'sd1189, 12'sd1865}, {12'sd-1169, 12'sd1490, 6'sd16}},
{{12'sd1989, 12'sd-1823, 13'sd2310}, {13'sd2077, 13'sd-2184, 12'sd1080}, {10'sd-324, 8'sd-103, 13'sd2079}},
{{11'sd-584, 11'sd-739, 13'sd-2056}, {11'sd831, 11'sd730, 12'sd-1646}, {10'sd316, 11'sd-568, 10'sd446}},
{{12'sd2039, 11'sd533, 10'sd358}, {12'sd1535, 10'sd274, 12'sd-1413}, {13'sd-2064, 13'sd-2763, 13'sd2203}},
{{12'sd1289, 9'sd158, 10'sd316}, {12'sd1215, 10'sd506, 9'sd209}, {9'sd-138, 11'sd-766, 12'sd1346}},
{{13'sd-2413, 12'sd-1761, 5'sd-8}, {13'sd3203, 12'sd-1049, 12'sd1065}, {11'sd881, 12'sd2042, 11'sd-720}},
{{13'sd-3103, 12'sd1938, 12'sd1268}, {13'sd2329, 12'sd1888, 12'sd-1472}, {13'sd2106, 12'sd-1584, 12'sd1043}}},
{
{{12'sd-1316, 12'sd-1535, 12'sd1257}, {12'sd1242, 13'sd-2960, 12'sd-1239}, {11'sd844, 12'sd-1658, 12'sd1683}},
{{12'sd1721, 12'sd1289, 12'sd-1889}, {12'sd1699, 13'sd-2371, 9'sd-138}, {12'sd1718, 12'sd-1670, 12'sd-1817}},
{{12'sd-1381, 12'sd1918, 13'sd-2413}, {11'sd952, 9'sd244, 11'sd-995}, {12'sd1537, 12'sd1278, 12'sd-1529}},
{{12'sd-1734, 12'sd-1527, 12'sd-1335}, {10'sd286, 10'sd-321, 12'sd1425}, {11'sd802, 12'sd-1792, 13'sd3635}},
{{12'sd1538, 9'sd-189, 13'sd2385}, {11'sd1023, 13'sd-3667, 13'sd-2172}, {11'sd-740, 14'sd-6018, 14'sd-6010}},
{{13'sd3487, 14'sd-5131, 10'sd-354}, {14'sd4660, 13'sd-2491, 5'sd-9}, {13'sd2693, 12'sd-1247, 12'sd-1587}},
{{13'sd2237, 14'sd-6487, 15'sd-8205}, {13'sd3167, 13'sd-2840, 14'sd-6078}, {14'sd5699, 13'sd-2230, 11'sd856}},
{{11'sd850, 13'sd-2804, 12'sd1809}, {11'sd-566, 13'sd-3066, 9'sd-133}, {13'sd-2122, 11'sd926, 12'sd-1846}},
{{9'sd159, 9'sd178, 11'sd-763}, {13'sd2735, 9'sd159, 12'sd1572}, {12'sd1192, 12'sd-1996, 11'sd-884}},
{{11'sd920, 10'sd442, 12'sd1617}, {13'sd3017, 12'sd-1651, 13'sd-2478}, {11'sd-787, 13'sd2180, 12'sd-1609}},
{{12'sd1536, 11'sd793, 11'sd-720}, {10'sd361, 13'sd2443, 10'sd494}, {12'sd1397, 13'sd2153, 12'sd-1275}},
{{8'sd74, 12'sd1034, 13'sd4010}, {11'sd-741, 11'sd536, 8'sd94}, {10'sd436, 13'sd-2102, 12'sd1134}},
{{13'sd3293, 11'sd583, 12'sd-2014}, {10'sd-447, 10'sd369, 13'sd-3625}, {12'sd-1183, 11'sd950, 12'sd1125}},
{{9'sd-254, 10'sd-509, 12'sd1273}, {12'sd1549, 13'sd2655, 12'sd1116}, {13'sd-2450, 13'sd-2549, 9'sd-136}},
{{13'sd2906, 15'sd8857, 13'sd3030}, {14'sd6725, 13'sd3691, 13'sd3454}, {11'sd902, 14'sd4146, 11'sd911}},
{{12'sd-1890, 12'sd1195, 13'sd3334}, {11'sd856, 12'sd-1366, 11'sd758}, {10'sd442, 12'sd-1866, 12'sd1754}},
{{12'sd1897, 12'sd-1113, 12'sd1095}, {13'sd-3190, 12'sd1431, 10'sd-438}, {11'sd-590, 12'sd1056, 10'sd-368}},
{{14'sd5927, 13'sd4091, 11'sd942}, {13'sd2416, 11'sd976, 11'sd-969}, {13'sd2260, 13'sd2260, 9'sd-233}},
{{12'sd-1411, 11'sd-676, 10'sd-468}, {13'sd3030, 10'sd344, 13'sd2067}, {13'sd2073, 10'sd342, 10'sd495}},
{{12'sd-1484, 11'sd-582, 12'sd-1217}, {12'sd-1221, 12'sd-1526, 12'sd-1696}, {12'sd-1329, 8'sd110, 13'sd2534}},
{{13'sd-3347, 12'sd-1051, 13'sd-2995}, {8'sd-97, 12'sd1443, 13'sd-2698}, {9'sd-215, 12'sd1314, 9'sd-150}},
{{9'sd228, 5'sd12, 11'sd575}, {11'sd1019, 10'sd260, 12'sd1201}, {11'sd830, 12'sd1444, 13'sd2304}},
{{12'sd1638, 12'sd-1246, 12'sd2041}, {12'sd1508, 12'sd-1883, 11'sd914}, {12'sd-1155, 11'sd978, 12'sd1680}},
{{13'sd-2563, 13'sd2383, 8'sd-127}, {12'sd1766, 13'sd2459, 12'sd-1112}, {10'sd-453, 10'sd-422, 12'sd1382}},
{{12'sd-1045, 12'sd-1983, 10'sd308}, {4'sd7, 13'sd-2613, 9'sd-150}, {12'sd-1265, 11'sd1017, 11'sd846}},
{{13'sd2689, 13'sd2590, 12'sd1893}, {10'sd-459, 13'sd-2365, 12'sd1740}, {12'sd1548, 12'sd1176, 13'sd-2439}},
{{13'sd-2550, 12'sd-1356, 12'sd-1734}, {12'sd-1043, 12'sd-1457, 13'sd-3394}, {11'sd618, 9'sd212, 13'sd-3951}},
{{11'sd714, 12'sd1705, 12'sd1460}, {13'sd2352, 13'sd-2133, 8'sd-70}, {12'sd1699, 13'sd2116, 12'sd1522}},
{{12'sd1249, 12'sd1462, 10'sd-328}, {12'sd1545, 13'sd3591, 12'sd1870}, {9'sd-230, 10'sd503, 10'sd260}},
{{10'sd470, 13'sd-2840, 10'sd496}, {12'sd1457, 12'sd1315, 12'sd1753}, {12'sd-1063, 11'sd-655, 12'sd1125}},
{{12'sd-1534, 13'sd2367, 11'sd-685}, {13'sd2073, 13'sd-2813, 11'sd612}, {10'sd292, 12'sd1419, 12'sd-1602}},
{{13'sd-3373, 13'sd2586, 12'sd1814}, {11'sd-743, 12'sd1408, 13'sd2888}, {12'sd1474, 10'sd427, 12'sd-1483}},
{{11'sd691, 12'sd1125, 13'sd2102}, {13'sd-3400, 13'sd-2120, 13'sd2719}, {13'sd-3169, 12'sd1924, 12'sd1261}},
{{12'sd-1217, 13'sd3105, 13'sd2266}, {10'sd-271, 11'sd-737, 9'sd247}, {9'sd-162, 14'sd4346, 13'sd3069}},
{{9'sd-195, 13'sd2563, 9'sd-141}, {13'sd-2792, 13'sd-2321, 11'sd-744}, {11'sd-921, 10'sd353, 12'sd1170}},
{{9'sd-155, 13'sd-2116, 12'sd1531}, {11'sd586, 10'sd473, 10'sd-353}, {10'sd376, 10'sd486, 12'sd1269}},
{{14'sd-7923, 9'sd-147, 12'sd-1793}, {14'sd-4103, 13'sd2215, 11'sd716}, {12'sd-1673, 13'sd2210, 12'sd1601}},
{{10'sd459, 11'sd-865, 12'sd1195}, {12'sd1603, 12'sd1241, 13'sd-3013}, {13'sd3863, 13'sd2505, 12'sd-1869}},
{{12'sd-1804, 12'sd-1213, 11'sd-772}, {12'sd1333, 13'sd2352, 11'sd-719}, {13'sd-3020, 13'sd-2192, 13'sd-2198}},
{{13'sd2936, 12'sd1831, 12'sd-1211}, {13'sd-2064, 12'sd-1649, 10'sd-375}, {10'sd474, 12'sd-1827, 13'sd-2992}},
{{12'sd1229, 12'sd-2011, 13'sd-2589}, {11'sd-1012, 11'sd786, 9'sd158}, {11'sd961, 6'sd24, 11'sd-1016}},
{{11'sd668, 13'sd3044, 12'sd1833}, {12'sd1636, 9'sd129, 12'sd-1371}, {12'sd-1036, 13'sd-2912, 14'sd-4700}},
{{11'sd515, 11'sd-960, 11'sd-1021}, {11'sd789, 13'sd2066, 13'sd-3090}, {14'sd5840, 14'sd4841, 11'sd-567}},
{{13'sd-2618, 13'sd-2243, 14'sd-5771}, {14'sd-4912, 14'sd-6093, 14'sd-5242}, {14'sd-7801, 13'sd-3810, 15'sd-11710}},
{{11'sd619, 13'sd2200, 12'sd-1191}, {12'sd1741, 11'sd-983, 11'sd-928}, {11'sd740, 11'sd565, 12'sd-1561}},
{{13'sd-3196, 12'sd1263, 11'sd-656}, {12'sd-1177, 11'sd702, 11'sd1002}, {10'sd-508, 10'sd416, 13'sd2267}},
{{13'sd-3995, 13'sd2108, 13'sd2360}, {8'sd73, 12'sd1328, 13'sd3208}, {11'sd611, 12'sd1871, 14'sd5536}},
{{12'sd-1335, 12'sd1072, 11'sd-1014}, {11'sd-835, 11'sd769, 13'sd-2168}, {11'sd862, 12'sd1130, 11'sd-530}},
{{10'sd448, 12'sd-1789, 13'sd-2857}, {12'sd1334, 10'sd-392, 10'sd-356}, {9'sd207, 13'sd3726, 13'sd2921}},
{{14'sd-4401, 11'sd850, 12'sd1242}, {13'sd-2753, 9'sd-203, 13'sd3440}, {14'sd-5245, 13'sd-2852, 11'sd753}},
{{10'sd-322, 13'sd3749, 12'sd1444}, {8'sd-94, 12'sd1038, 12'sd1508}, {12'sd-1320, 13'sd2817, 12'sd1041}},
{{11'sd689, 11'sd870, 11'sd644}, {12'sd1680, 9'sd-172, 8'sd73}, {13'sd2077, 13'sd-3567, 12'sd1488}},
{{12'sd1457, 12'sd1252, 11'sd1006}, {13'sd2607, 13'sd-2311, 12'sd-1037}, {10'sd-401, 13'sd-3026, 13'sd-3390}},
{{11'sd836, 13'sd-3042, 13'sd-2568}, {10'sd384, 13'sd-2116, 12'sd1129}, {13'sd3228, 13'sd2061, 11'sd831}},
{{11'sd826, 13'sd-2379, 14'sd-4588}, {5'sd11, 13'sd2208, 14'sd-4580}, {10'sd467, 13'sd2743, 10'sd-326}},
{{13'sd-3710, 13'sd-3510, 12'sd1089}, {12'sd-1714, 12'sd1275, 12'sd-1305}, {13'sd-3408, 13'sd2204, 12'sd1977}},
{{13'sd-2065, 12'sd-1773, 13'sd-2384}, {13'sd-3734, 10'sd462, 13'sd-3054}, {14'sd-5321, 14'sd-5891, 14'sd-5559}},
{{13'sd2254, 11'sd971, 13'sd2213}, {14'sd4571, 13'sd3142, 11'sd-797}, {12'sd1861, 11'sd-836, 12'sd-1874}},
{{13'sd2309, 9'sd252, 13'sd-2244}, {13'sd2701, 11'sd1022, 13'sd-3176}, {12'sd1299, 13'sd-2072, 12'sd-1818}},
{{11'sd590, 11'sd654, 11'sd955}, {10'sd-337, 13'sd3019, 12'sd1109}, {15'sd13292, 14'sd6569, 15'sd8743}},
{{12'sd-2034, 11'sd-587, 10'sd293}, {13'sd-3048, 12'sd1758, 11'sd-513}, {9'sd-174, 13'sd2260, 8'sd-71}},
{{11'sd-536, 11'sd-670, 13'sd2790}, {11'sd824, 13'sd-2356, 12'sd1047}, {11'sd985, 13'sd-2757, 11'sd-697}},
{{13'sd-2841, 12'sd-1656, 10'sd-435}, {13'sd-3441, 11'sd-892, 7'sd50}, {12'sd-1349, 14'sd-4740, 12'sd1852}},
{{11'sd-597, 11'sd561, 10'sd373}, {12'sd1806, 10'sd-329, 9'sd161}, {13'sd2683, 13'sd2255, 13'sd2388}}},
{
{{10'sd511, 13'sd-2731, 12'sd-1676}, {12'sd-1577, 11'sd1017, 8'sd69}, {11'sd833, 12'sd1136, 13'sd2768}},
{{11'sd571, 12'sd-2044, 12'sd-1685}, {6'sd-31, 10'sd-385, 12'sd-1340}, {12'sd1559, 10'sd-358, 12'sd-1751}},
{{12'sd-1594, 11'sd886, 13'sd2134}, {13'sd2576, 9'sd147, 12'sd-1418}, {12'sd1624, 13'sd-2105, 11'sd720}},
{{10'sd483, 13'sd2289, 9'sd233}, {12'sd-1644, 12'sd1677, 12'sd1828}, {13'sd2864, 11'sd-724, 12'sd-1395}},
{{13'sd3615, 12'sd1961, 12'sd1623}, {13'sd2615, 10'sd461, 13'sd2972}, {11'sd611, 13'sd-2107, 11'sd726}},
{{9'sd172, 8'sd96, 13'sd-3316}, {12'sd-1661, 12'sd-1829, 10'sd-321}, {13'sd-2800, 12'sd1560, 13'sd2185}},
{{13'sd-2664, 12'sd1543, 12'sd1954}, {12'sd1773, 13'sd2457, 12'sd1266}, {8'sd108, 13'sd2121, 13'sd2652}},
{{12'sd-1595, 11'sd824, 9'sd160}, {12'sd-1423, 12'sd1728, 7'sd36}, {12'sd-1353, 11'sd849, 12'sd-1040}},
{{12'sd-1405, 13'sd-2557, 9'sd209}, {11'sd-770, 12'sd1548, 13'sd-2144}, {12'sd-1540, 13'sd2179, 12'sd1043}},
{{13'sd-2149, 10'sd-457, 13'sd2112}, {8'sd104, 13'sd2413, 13'sd-2146}, {12'sd-1051, 11'sd757, 13'sd2143}},
{{12'sd1996, 10'sd502, 12'sd1417}, {8'sd-126, 9'sd-166, 13'sd2753}, {10'sd-480, 12'sd-2005, 9'sd235}},
{{13'sd2366, 13'sd-2155, 13'sd2578}, {6'sd22, 13'sd-2942, 12'sd-1504}, {12'sd-1905, 13'sd-2663, 13'sd-2287}},
{{12'sd-1529, 11'sd929, 12'sd1043}, {13'sd-2219, 12'sd1151, 12'sd-1712}, {9'sd-169, 10'sd-392, 12'sd1280}},
{{12'sd-1665, 12'sd1161, 12'sd-1607}, {13'sd-2122, 13'sd2233, 10'sd398}, {12'sd-1878, 13'sd-2339, 11'sd-953}},
{{10'sd-314, 12'sd-1457, 13'sd2048}, {11'sd-655, 12'sd-1637, 12'sd1567}, {12'sd1687, 11'sd-929, 12'sd-1451}},
{{12'sd1786, 9'sd210, 11'sd656}, {11'sd778, 11'sd869, 11'sd904}, {13'sd2557, 13'sd2582, 11'sd659}},
{{11'sd-756, 12'sd-1972, 13'sd-2511}, {12'sd1207, 10'sd356, 11'sd597}, {13'sd2735, 12'sd-1398, 13'sd-2680}},
{{12'sd-1623, 12'sd1235, 11'sd666}, {12'sd-1192, 13'sd2375, 13'sd2341}, {11'sd-710, 12'sd-1922, 12'sd1202}},
{{11'sd-870, 12'sd1210, 11'sd-690}, {12'sd1164, 13'sd-2133, 8'sd70}, {13'sd-2210, 12'sd-1923, 12'sd-1238}},
{{12'sd1690, 8'sd74, 12'sd-1798}, {13'sd2870, 12'sd-1246, 12'sd1379}, {11'sd534, 11'sd981, 11'sd786}},
{{12'sd1786, 11'sd-769, 12'sd-1707}, {12'sd1281, 12'sd-1177, 11'sd734}, {13'sd-2221, 13'sd2957, 12'sd-1199}},
{{12'sd-1801, 12'sd-1232, 12'sd1637}, {12'sd2006, 10'sd327, 10'sd463}, {12'sd1377, 10'sd-359, 12'sd-1079}},
{{11'sd919, 12'sd1962, 10'sd433}, {12'sd-1652, 9'sd130, 13'sd-2130}, {12'sd1787, 12'sd-1571, 13'sd-2569}},
{{9'sd155, 13'sd-2353, 9'sd165}, {13'sd2735, 12'sd-1869, 11'sd-692}, {12'sd-1749, 10'sd344, 12'sd-1202}},
{{7'sd54, 13'sd2915, 8'sd-102}, {13'sd-2190, 13'sd-2129, 13'sd-2211}, {12'sd-1632, 13'sd2108, 13'sd2713}},
{{7'sd40, 12'sd-1477, 10'sd-338}, {12'sd-1316, 13'sd-2439, 13'sd2248}, {11'sd644, 13'sd2570, 11'sd-664}},
{{12'sd-1144, 13'sd2241, 12'sd1032}, {14'sd4822, 14'sd4910, 9'sd142}, {13'sd2558, 14'sd4252, 13'sd3356}},
{{11'sd689, 12'sd1797, 13'sd2066}, {13'sd2557, 8'sd-110, 11'sd641}, {12'sd-1278, 8'sd91, 6'sd16}},
{{12'sd-1027, 10'sd323, 13'sd3519}, {11'sd997, 13'sd-2305, 13'sd2359}, {11'sd-770, 13'sd-2649, 13'sd2463}},
{{11'sd-927, 9'sd255, 12'sd-1629}, {12'sd1777, 11'sd956, 11'sd-832}, {12'sd-1547, 12'sd1220, 13'sd2639}},
{{12'sd-1563, 13'sd-2196, 13'sd-2646}, {12'sd-1522, 13'sd2305, 12'sd-1505}, {10'sd-344, 12'sd-1805, 11'sd760}},
{{11'sd-763, 13'sd-2266, 12'sd1519}, {13'sd-2896, 11'sd-815, 1'sd0}, {12'sd2015, 12'sd-1750, 11'sd639}},
{{12'sd1390, 9'sd151, 12'sd-1600}, {12'sd-1085, 13'sd2457, 12'sd-1178}, {12'sd-1832, 9'sd250, 11'sd-996}},
{{12'sd1156, 12'sd1742, 13'sd2357}, {7'sd59, 11'sd914, 12'sd1734}, {11'sd1007, 10'sd488, 12'sd1392}},
{{9'sd154, 10'sd-508, 13'sd-2707}, {12'sd-1990, 10'sd424, 10'sd360}, {11'sd-588, 13'sd-2582, 13'sd-2637}},
{{10'sd264, 11'sd-565, 11'sd-870}, {12'sd1718, 12'sd1816, 13'sd2499}, {12'sd-1473, 9'sd172, 12'sd-2036}},
{{12'sd-1620, 11'sd-996, 11'sd-598}, {13'sd2712, 11'sd1008, 13'sd-2072}, {10'sd-432, 12'sd-2010, 12'sd-1913}},
{{12'sd-1029, 13'sd2075, 13'sd-2352}, {12'sd-1752, 11'sd-560, 12'sd1399}, {12'sd1913, 11'sd-610, 10'sd502}},
{{9'sd-141, 11'sd-800, 13'sd-2537}, {12'sd1778, 12'sd1843, 13'sd2643}, {11'sd-659, 12'sd1267, 12'sd1449}},
{{13'sd-2268, 12'sd-2022, 10'sd303}, {9'sd-217, 13'sd2101, 4'sd4}, {11'sd-546, 12'sd-1752, 12'sd1575}},
{{12'sd-1279, 13'sd2346, 12'sd-1620}, {13'sd2061, 13'sd2125, 12'sd1511}, {11'sd764, 13'sd2716, 12'sd1062}},
{{10'sd445, 11'sd-875, 12'sd1460}, {6'sd-31, 12'sd-1607, 10'sd-382}, {12'sd1783, 10'sd397, 12'sd-1188}},
{{13'sd2986, 13'sd2117, 12'sd1647}, {7'sd-61, 11'sd574, 13'sd3161}, {13'sd2286, 11'sd-613, 12'sd-1652}},
{{12'sd1225, 10'sd396, 12'sd1197}, {12'sd1360, 13'sd3381, 12'sd1826}, {12'sd-1802, 8'sd91, 12'sd1999}},
{{13'sd-2178, 9'sd-178, 13'sd2203}, {12'sd-1408, 12'sd1852, 12'sd1109}, {13'sd-2693, 13'sd-2535, 13'sd-2423}},
{{9'sd132, 13'sd2716, 12'sd1990}, {11'sd574, 12'sd1677, 10'sd-365}, {12'sd-1817, 12'sd1239, 8'sd-72}},
{{13'sd-2625, 13'sd2218, 10'sd-367}, {12'sd1502, 11'sd-769, 13'sd-2155}, {12'sd-1395, 13'sd2746, 6'sd26}},
{{12'sd1994, 13'sd3561, 10'sd-426}, {11'sd-941, 12'sd-1049, 10'sd330}, {13'sd2703, 11'sd-978, 12'sd1633}},
{{13'sd2721, 13'sd-2306, 10'sd-271}, {12'sd1776, 12'sd1663, 13'sd-2344}, {12'sd1378, 13'sd2372, 12'sd-1794}},
{{13'sd-2161, 10'sd-429, 12'sd-1697}, {13'sd-2389, 13'sd-2346, 13'sd-3003}, {11'sd600, 9'sd-223, 11'sd-861}},
{{11'sd819, 8'sd-88, 12'sd1293}, {12'sd-1991, 12'sd-1776, 12'sd1972}, {10'sd-295, 13'sd-2143, 12'sd-1582}},
{{11'sd-709, 10'sd-279, 12'sd1178}, {13'sd-2533, 12'sd1799, 12'sd-1878}, {10'sd323, 11'sd-738, 12'sd-1578}},
{{10'sd-341, 11'sd-849, 8'sd121}, {7'sd46, 12'sd-1637, 12'sd1111}, {12'sd-1708, 13'sd-2412, 13'sd2088}},
{{11'sd932, 13'sd2644, 10'sd-404}, {12'sd1451, 12'sd1385, 12'sd1764}, {12'sd1988, 13'sd2977, 12'sd1759}},
{{12'sd-1149, 11'sd863, 12'sd-1184}, {12'sd1689, 13'sd2205, 12'sd1249}, {13'sd2554, 12'sd1836, 11'sd857}},
{{11'sd608, 12'sd-1865, 11'sd-824}, {7'sd49, 9'sd-188, 3'sd2}, {12'sd1841, 12'sd1118, 12'sd1506}},
{{13'sd-2669, 12'sd1725, 13'sd-2061}, {12'sd-1806, 11'sd965, 13'sd-2172}, {10'sd-391, 12'sd1278, 12'sd1298}},
{{12'sd-1750, 10'sd-404, 10'sd-390}, {12'sd-2012, 12'sd1845, 13'sd2484}, {13'sd2299, 10'sd416, 13'sd-3303}},
{{13'sd2608, 12'sd2036, 8'sd-80}, {11'sd-831, 13'sd-2222, 9'sd179}, {13'sd-2355, 11'sd980, 12'sd1221}},
{{13'sd3723, 8'sd-122, 13'sd3176}, {12'sd-1354, 11'sd-762, 13'sd3238}, {13'sd-2207, 11'sd-949, 13'sd2469}},
{{13'sd2871, 9'sd239, 12'sd-1339}, {13'sd2271, 13'sd-2740, 13'sd2119}, {11'sd564, 13'sd-2317, 12'sd-1781}},
{{12'sd1746, 12'sd1500, 10'sd-352}, {12'sd1237, 11'sd582, 13'sd2578}, {12'sd-1585, 10'sd365, 12'sd1194}},
{{5'sd8, 11'sd794, 12'sd-1971}, {12'sd-1737, 10'sd344, 13'sd2097}, {9'sd-187, 11'sd611, 11'sd-525}},
{{12'sd1285, 13'sd-2367, 11'sd-753}, {10'sd-487, 12'sd-1472, 12'sd1456}, {9'sd-133, 11'sd581, 8'sd91}}},
{
{{12'sd-1467, 12'sd-1565, 9'sd185}, {12'sd-1313, 11'sd991, 9'sd171}, {12'sd1690, 11'sd-999, 12'sd1636}},
{{11'sd694, 13'sd2572, 9'sd164}, {13'sd2490, 10'sd396, 12'sd1614}, {12'sd1749, 13'sd-2133, 12'sd1396}},
{{13'sd2796, 7'sd-33, 12'sd1225}, {11'sd759, 13'sd-2200, 8'sd-110}, {12'sd1765, 12'sd-1943, 11'sd689}},
{{12'sd1041, 11'sd720, 13'sd2356}, {13'sd2448, 12'sd1872, 11'sd-798}, {12'sd-1191, 13'sd-2351, 12'sd-1160}},
{{10'sd303, 11'sd-977, 12'sd1550}, {11'sd712, 7'sd-55, 13'sd-3406}, {10'sd-414, 13'sd-3539, 12'sd-1752}},
{{13'sd-2914, 13'sd2304, 10'sd-412}, {10'sd-386, 13'sd2923, 12'sd-1290}, {12'sd-1452, 10'sd275, 13'sd3367}},
{{12'sd-2040, 12'sd1529, 10'sd457}, {11'sd-640, 11'sd531, 11'sd905}, {12'sd-1188, 13'sd2245, 10'sd-298}},
{{13'sd2628, 13'sd2250, 13'sd-2615}, {12'sd1226, 12'sd1195, 9'sd-241}, {12'sd-1811, 11'sd645, 13'sd2130}},
{{12'sd1361, 13'sd-2139, 13'sd2115}, {12'sd-1782, 12'sd1804, 13'sd2338}, {13'sd-2874, 11'sd519, 10'sd-297}},
{{13'sd-2173, 11'sd-995, 13'sd2351}, {12'sd1394, 12'sd1565, 12'sd-1649}, {13'sd-2332, 12'sd1175, 8'sd106}},
{{13'sd2561, 13'sd2281, 12'sd-1509}, {12'sd1174, 13'sd2402, 10'sd328}, {9'sd239, 11'sd-865, 7'sd51}},
{{12'sd-1170, 9'sd-239, 12'sd-1359}, {12'sd1323, 11'sd-915, 9'sd-223}, {10'sd273, 12'sd1562, 11'sd-552}},
{{6'sd31, 12'sd-1203, 13'sd-2888}, {9'sd162, 13'sd-3035, 13'sd-3668}, {13'sd-2593, 11'sd-647, 12'sd-1217}},
{{12'sd-1703, 11'sd702, 13'sd-2503}, {12'sd1177, 12'sd-1095, 12'sd-1643}, {12'sd-1084, 9'sd-234, 12'sd-1377}},
{{13'sd2874, 12'sd1725, 10'sd363}, {12'sd1631, 11'sd-798, 11'sd966}, {12'sd-1160, 10'sd-315, 11'sd601}},
{{12'sd1602, 10'sd511, 9'sd231}, {13'sd2528, 12'sd-1031, 11'sd-789}, {12'sd-1178, 12'sd1063, 13'sd-2164}},
{{10'sd-371, 13'sd-2478, 12'sd-1600}, {11'sd992, 11'sd-884, 13'sd-2337}, {13'sd2795, 12'sd1598, 8'sd67}},
{{5'sd-10, 7'sd42, 12'sd-1283}, {10'sd-504, 11'sd982, 12'sd-1619}, {13'sd-2305, 12'sd1921, 11'sd1004}},
{{12'sd1158, 10'sd277, 12'sd-1846}, {13'sd-2288, 8'sd-71, 12'sd1059}, {12'sd1873, 11'sd-674, 11'sd790}},
{{10'sd325, 9'sd136, 12'sd-1320}, {13'sd2540, 12'sd-1281, 13'sd-2384}, {12'sd1812, 11'sd-860, 13'sd-2226}},
{{12'sd-2039, 12'sd-1105, 12'sd1704}, {12'sd-1475, 12'sd1949, 11'sd902}, {10'sd301, 8'sd-65, 13'sd-2218}},
{{13'sd2097, 11'sd630, 12'sd-1045}, {12'sd1487, 13'sd2176, 13'sd2502}, {12'sd-1101, 11'sd527, 11'sd742}},
{{12'sd1317, 12'sd-1248, 13'sd-2773}, {13'sd-2514, 9'sd-150, 13'sd-2337}, {13'sd2325, 9'sd-252, 11'sd556}},
{{11'sd872, 13'sd2237, 13'sd-2434}, {11'sd680, 12'sd1601, 12'sd-1532}, {13'sd-2611, 10'sd466, 13'sd-2320}},
{{12'sd1500, 8'sd65, 12'sd-1400}, {13'sd-2433, 12'sd1838, 12'sd-1045}, {12'sd1406, 9'sd-181, 12'sd-1178}},
{{13'sd-2249, 12'sd1687, 11'sd-618}, {11'sd692, 13'sd-2351, 12'sd1394}, {13'sd2445, 11'sd-849, 12'sd-1479}},
{{12'sd-1193, 13'sd2068, 11'sd609}, {11'sd1008, 12'sd1077, 13'sd2918}, {13'sd2309, 12'sd-1949, 13'sd2348}},
{{12'sd-1530, 13'sd-2192, 11'sd628}, {9'sd-217, 7'sd55, 12'sd-1765}, {11'sd-745, 12'sd-1400, 13'sd-2529}},
{{12'sd-1451, 13'sd-2397, 12'sd1221}, {12'sd1824, 13'sd2460, 13'sd-2255}, {11'sd838, 13'sd-2429, 12'sd-1752}},
{{11'sd-904, 9'sd200, 12'sd1340}, {13'sd-2562, 12'sd1485, 13'sd-2528}, {12'sd-1211, 9'sd229, 12'sd-1252}},
{{12'sd-1858, 12'sd1967, 12'sd-1989}, {11'sd543, 13'sd2444, 12'sd1131}, {11'sd-633, 11'sd554, 13'sd-2511}},
{{10'sd496, 12'sd-1283, 13'sd2761}, {12'sd-1203, 10'sd411, 12'sd-1816}, {13'sd-2072, 13'sd2223, 13'sd-2410}},
{{11'sd607, 6'sd24, 11'sd772}, {13'sd-2629, 12'sd1557, 12'sd-1225}, {12'sd1606, 13'sd-2128, 11'sd821}},
{{12'sd1148, 12'sd-1403, 12'sd-1400}, {11'sd-1018, 12'sd1654, 11'sd-997}, {12'sd1718, 13'sd-2241, 10'sd-407}},
{{10'sd302, 13'sd2154, 12'sd-1469}, {12'sd-1502, 12'sd-1440, 11'sd-895}, {11'sd705, 12'sd1691, 13'sd2449}},
{{13'sd-2312, 12'sd1665, 12'sd-1844}, {12'sd1102, 12'sd1756, 13'sd2452}, {10'sd-367, 13'sd-2199, 9'sd196}},
{{12'sd-1898, 9'sd-219, 12'sd-1482}, {13'sd-2409, 13'sd2267, 13'sd3098}, {9'sd-242, 10'sd-310, 13'sd2544}},
{{12'sd1604, 13'sd-2694, 12'sd1581}, {12'sd1042, 13'sd-2962, 11'sd525}, {11'sd-696, 13'sd-2474, 11'sd-650}},
{{10'sd281, 13'sd-2357, 12'sd1451}, {13'sd2393, 12'sd1118, 9'sd-229}, {13'sd2485, 13'sd2699, 13'sd2570}},
{{13'sd-2301, 12'sd1226, 8'sd-108}, {12'sd-1394, 12'sd-1929, 6'sd-23}, {12'sd1350, 13'sd-2456, 11'sd721}},
{{9'sd130, 13'sd-2308, 11'sd810}, {12'sd-1049, 11'sd-519, 11'sd972}, {9'sd-255, 12'sd-1625, 11'sd-772}},
{{13'sd-2067, 13'sd-2308, 11'sd785}, {12'sd-1859, 13'sd-2153, 13'sd-2822}, {12'sd-1798, 12'sd1524, 13'sd-2342}},
{{12'sd-1522, 11'sd-515, 11'sd-911}, {11'sd-928, 12'sd1272, 11'sd572}, {10'sd297, 12'sd-1930, 13'sd2071}},
{{12'sd1978, 10'sd274, 13'sd2958}, {11'sd-668, 12'sd1957, 12'sd-1821}, {13'sd2306, 12'sd-1974, 12'sd1105}},
{{11'sd-881, 12'sd1955, 8'sd-123}, {12'sd-1657, 11'sd-593, 11'sd639}, {11'sd-590, 12'sd1639, 12'sd1171}},
{{11'sd884, 12'sd1999, 13'sd2439}, {7'sd-33, 12'sd1116, 13'sd-2181}, {12'sd1074, 12'sd2021, 12'sd-1958}},
{{12'sd1670, 13'sd-2475, 13'sd-3142}, {10'sd331, 11'sd695, 11'sd-686}, {11'sd726, 11'sd672, 10'sd384}},
{{9'sd-188, 13'sd2746, 13'sd-2155}, {12'sd-1408, 10'sd493, 12'sd1407}, {11'sd-934, 8'sd112, 12'sd-1154}},
{{8'sd-79, 13'sd2859, 13'sd3006}, {11'sd-945, 13'sd2765, 12'sd-1107}, {11'sd-1022, 9'sd-134, 12'sd1656}},
{{12'sd1629, 11'sd-620, 11'sd853}, {8'sd116, 10'sd-266, 13'sd-2402}, {12'sd1771, 6'sd30, 10'sd-448}},
{{13'sd-2273, 13'sd-2118, 12'sd-1780}, {12'sd-1703, 12'sd-1213, 11'sd-655}, {12'sd1201, 13'sd-2637, 10'sd380}},
{{12'sd1623, 11'sd-996, 9'sd-212}, {9'sd190, 10'sd273, 13'sd2100}, {12'sd-1661, 11'sd569, 13'sd-2485}},
{{12'sd-1376, 13'sd2646, 12'sd1473}, {12'sd1354, 12'sd-1612, 12'sd1401}, {11'sd538, 9'sd-242, 13'sd2156}},
{{8'sd-120, 12'sd1805, 13'sd2219}, {11'sd903, 12'sd-1315, 10'sd337}, {12'sd1070, 11'sd-572, 7'sd32}},
{{11'sd597, 13'sd-3065, 10'sd398}, {13'sd-3440, 11'sd884, 13'sd-2752}, {9'sd224, 8'sd74, 12'sd1597}},
{{9'sd-142, 13'sd-2095, 13'sd2662}, {12'sd-1213, 12'sd-1389, 11'sd-769}, {12'sd2019, 12'sd-1598, 12'sd-1842}},
{{11'sd-934, 13'sd-2641, 11'sd-610}, {13'sd-2312, 14'sd-4190, 14'sd-5680}, {13'sd-2238, 12'sd1035, 12'sd-1619}},
{{11'sd-601, 12'sd-1758, 12'sd1600}, {12'sd-1265, 11'sd-578, 13'sd-2728}, {11'sd-776, 8'sd84, 11'sd-774}},
{{13'sd2301, 12'sd-1284, 11'sd-920}, {11'sd-888, 11'sd-625, 12'sd-1085}, {12'sd1829, 13'sd2521, 13'sd-2154}},
{{10'sd-378, 13'sd2491, 13'sd2270}, {12'sd-1572, 10'sd508, 12'sd1114}, {12'sd-1989, 3'sd3, 8'sd106}},
{{12'sd-2011, 12'sd-1722, 12'sd1636}, {13'sd2089, 12'sd1143, 12'sd1198}, {10'sd423, 13'sd2607, 10'sd-260}},
{{10'sd-498, 11'sd-842, 10'sd-487}, {13'sd2484, 13'sd2058, 12'sd-1732}, {12'sd-1732, 12'sd-1736, 11'sd792}},
{{10'sd502, 10'sd344, 12'sd1778}, {13'sd-2212, 13'sd3047, 13'sd-2487}, {13'sd2157, 13'sd2775, 7'sd-43}},
{{11'sd-701, 12'sd1223, 12'sd-1459}, {13'sd2343, 11'sd666, 10'sd266}, {12'sd-1657, 12'sd-1158, 13'sd3114}}},
{
{{13'sd2657, 11'sd1020, 13'sd-2365}, {13'sd2521, 13'sd-2388, 12'sd1111}, {8'sd66, 12'sd-1903, 12'sd1966}},
{{13'sd2651, 13'sd2349, 11'sd974}, {12'sd2015, 13'sd2778, 13'sd-2086}, {12'sd2031, 11'sd752, 12'sd-1213}},
{{13'sd-2241, 11'sd661, 11'sd-693}, {13'sd-3128, 4'sd-7, 11'sd588}, {12'sd-1839, 11'sd-664, 12'sd-1218}},
{{12'sd1031, 10'sd-483, 13'sd2716}, {13'sd-2874, 10'sd467, 12'sd-1109}, {9'sd128, 12'sd-1582, 13'sd-2106}},
{{11'sd640, 10'sd490, 12'sd1700}, {11'sd686, 12'sd1411, 12'sd1779}, {14'sd-4526, 10'sd-347, 12'sd-1124}},
{{13'sd2052, 10'sd-273, 13'sd-2533}, {12'sd-1942, 13'sd-2586, 12'sd1812}, {12'sd-1999, 11'sd-674, 13'sd3919}},
{{13'sd-2253, 11'sd-752, 13'sd2892}, {13'sd-2411, 13'sd-2119, 7'sd51}, {12'sd1740, 13'sd-3961, 12'sd-1155}},
{{13'sd-3097, 12'sd1130, 10'sd484}, {11'sd727, 13'sd2369, 13'sd2584}, {12'sd-1208, 13'sd2303, 8'sd92}},
{{12'sd1218, 12'sd-1884, 12'sd1909}, {13'sd2624, 10'sd429, 13'sd-2117}, {7'sd-39, 12'sd-1957, 11'sd900}},
{{13'sd-2603, 12'sd-1504, 11'sd978}, {13'sd-2639, 13'sd2300, 11'sd1000}, {12'sd1879, 12'sd-1350, 12'sd1906}},
{{10'sd323, 13'sd2403, 12'sd-1583}, {13'sd-2658, 12'sd1535, 11'sd829}, {13'sd-3244, 12'sd2008, 12'sd-1921}},
{{10'sd-412, 11'sd619, 12'sd-1808}, {11'sd-687, 12'sd-1119, 11'sd753}, {9'sd218, 12'sd-2020, 12'sd-1315}},
{{12'sd1907, 13'sd2147, 12'sd-1586}, {13'sd3040, 12'sd1392, 8'sd113}, {12'sd-1950, 12'sd1894, 10'sd-303}},
{{12'sd1590, 12'sd-1633, 12'sd-1715}, {13'sd2355, 11'sd-549, 10'sd270}, {11'sd-640, 12'sd-1168, 12'sd-1933}},
{{11'sd-907, 11'sd-599, 12'sd-1440}, {12'sd-1156, 11'sd-749, 12'sd2046}, {3'sd-3, 9'sd-228, 11'sd780}},
{{12'sd2013, 12'sd1241, 12'sd1620}, {11'sd-939, 12'sd1737, 9'sd-209}, {10'sd-427, 13'sd-2310, 13'sd2586}},
{{11'sd795, 13'sd2583, 11'sd900}, {13'sd2267, 12'sd1841, 10'sd419}, {11'sd-881, 13'sd-2293, 10'sd-501}},
{{11'sd696, 11'sd-789, 12'sd1896}, {10'sd306, 12'sd1084, 13'sd3695}, {11'sd664, 8'sd-124, 13'sd3123}},
{{13'sd-2352, 12'sd1251, 12'sd1735}, {12'sd1553, 12'sd-1065, 12'sd-1533}, {11'sd-573, 11'sd-579, 13'sd2125}},
{{10'sd276, 10'sd382, 12'sd-1607}, {10'sd-362, 11'sd-563, 9'sd-213}, {13'sd2573, 13'sd2763, 13'sd-2541}},
{{9'sd-191, 12'sd-1039, 9'sd248}, {12'sd1681, 11'sd582, 12'sd1168}, {13'sd-2096, 13'sd-2698, 10'sd397}},
{{12'sd1480, 11'sd-772, 12'sd1074}, {13'sd2340, 13'sd2629, 9'sd-171}, {13'sd2767, 9'sd150, 12'sd1529}},
{{13'sd2596, 11'sd578, 13'sd-2208}, {12'sd1946, 12'sd-1815, 10'sd401}, {11'sd-664, 10'sd-269, 10'sd-500}},
{{12'sd-1117, 12'sd-1472, 13'sd-2103}, {13'sd-2160, 13'sd2166, 2'sd1}, {7'sd-44, 12'sd-1571, 12'sd1730}},
{{12'sd1918, 12'sd-1336, 12'sd-1300}, {12'sd-2001, 11'sd528, 10'sd364}, {13'sd2056, 12'sd1312, 13'sd3088}},
{{11'sd532, 11'sd-905, 10'sd428}, {12'sd-1651, 12'sd-1358, 13'sd2760}, {13'sd-3318, 13'sd2292, 12'sd-1178}},
{{11'sd-727, 13'sd-2870, 13'sd-3343}, {13'sd-2875, 12'sd-1850, 12'sd1873}, {10'sd482, 12'sd1461, 13'sd2332}},
{{10'sd347, 9'sd241, 11'sd-541}, {12'sd1686, 10'sd-389, 12'sd-1566}, {13'sd-3399, 12'sd1255, 12'sd-1888}},
{{12'sd1695, 7'sd-55, 12'sd-1041}, {10'sd305, 11'sd698, 13'sd2394}, {13'sd-2059, 10'sd-494, 6'sd-21}},
{{9'sd140, 13'sd-2879, 12'sd1346}, {9'sd-209, 12'sd-2042, 12'sd-1303}, {10'sd-476, 7'sd47, 12'sd1299}},
{{13'sd2456, 10'sd455, 9'sd-143}, {12'sd-1633, 10'sd-288, 12'sd-1544}, {13'sd-2292, 10'sd427, 12'sd1412}},
{{12'sd-1365, 12'sd1227, 12'sd-1392}, {10'sd-462, 12'sd1619, 12'sd-1180}, {13'sd2439, 12'sd-1470, 13'sd-2694}},
{{5'sd-14, 13'sd-2616, 13'sd2069}, {13'sd2263, 13'sd-2891, 13'sd2253}, {12'sd1525, 10'sd472, 9'sd-240}},
{{12'sd1904, 11'sd551, 12'sd1793}, {12'sd1934, 5'sd-8, 12'sd1928}, {13'sd2911, 12'sd-1537, 11'sd-523}},
{{13'sd2284, 10'sd-506, 14'sd-4273}, {13'sd-2401, 12'sd1722, 9'sd-194}, {13'sd3155, 12'sd1155, 4'sd-7}},
{{12'sd1985, 12'sd-1227, 13'sd-2775}, {12'sd-1440, 13'sd2491, 12'sd-1916}, {12'sd1658, 9'sd220, 12'sd1208}},
{{7'sd-54, 13'sd-3484, 14'sd-4222}, {12'sd-1950, 12'sd-1592, 14'sd-5477}, {13'sd2905, 11'sd-935, 14'sd-4557}},
{{12'sd1336, 12'sd-2045, 12'sd-2034}, {13'sd2145, 12'sd-1625, 13'sd-2797}, {12'sd1862, 13'sd3191, 12'sd1434}},
{{13'sd2065, 12'sd-1391, 10'sd-471}, {12'sd1131, 13'sd-2742, 13'sd2363}, {12'sd-1863, 11'sd855, 12'sd-1886}},
{{12'sd-1241, 13'sd2341, 12'sd1387}, {12'sd1805, 12'sd1795, 10'sd-357}, {12'sd-1916, 12'sd1600, 12'sd-1551}},
{{13'sd-2220, 11'sd844, 11'sd637}, {12'sd-1587, 12'sd-1601, 11'sd839}, {11'sd-695, 13'sd2344, 12'sd1900}},
{{12'sd1320, 12'sd-1245, 11'sd-939}, {12'sd1161, 12'sd1417, 13'sd-3367}, {13'sd-2506, 13'sd-3524, 13'sd-2394}},
{{14'sd-4441, 12'sd-1249, 10'sd337}, {14'sd-4496, 13'sd-2558, 13'sd2700}, {11'sd-746, 13'sd-2650, 12'sd1038}},
{{12'sd-1970, 13'sd-3843, 11'sd-540}, {9'sd178, 12'sd1303, 10'sd-321}, {12'sd1736, 13'sd-3625, 14'sd-4741}},
{{11'sd584, 12'sd1865, 11'sd-645}, {13'sd2578, 12'sd1289, 12'sd2004}, {11'sd1018, 11'sd852, 10'sd-272}},
{{13'sd-2429, 12'sd-1848, 12'sd1542}, {9'sd-242, 12'sd-1671, 12'sd1515}, {13'sd2741, 12'sd-1058, 9'sd-136}},
{{9'sd-230, 9'sd149, 7'sd-61}, {10'sd-297, 13'sd-2364, 13'sd-2684}, {11'sd-921, 8'sd-74, 12'sd1237}},
{{11'sd-670, 12'sd-1735, 13'sd-2375}, {11'sd925, 13'sd-2138, 13'sd3123}, {10'sd435, 12'sd-1210, 13'sd-3264}},
{{13'sd-2849, 11'sd-932, 10'sd478}, {12'sd-1044, 12'sd-1423, 13'sd3039}, {11'sd-1017, 10'sd-359, 9'sd-137}},
{{13'sd3389, 8'sd78, 12'sd1279}, {13'sd2224, 13'sd2576, 12'sd1942}, {13'sd-2761, 13'sd-3063, 13'sd2549}},
{{12'sd1138, 10'sd-425, 13'sd-2929}, {13'sd3053, 12'sd-1364, 13'sd2206}, {12'sd1449, 9'sd-189, 12'sd-1630}},
{{12'sd-1858, 8'sd122, 11'sd-990}, {13'sd2281, 11'sd-651, 12'sd1098}, {11'sd786, 12'sd-1317, 12'sd-1138}},
{{12'sd1990, 12'sd1130, 10'sd-261}, {12'sd1081, 11'sd588, 11'sd-784}, {13'sd-3685, 14'sd-5105, 10'sd-497}},
{{11'sd-690, 12'sd1850, 12'sd1186}, {11'sd556, 12'sd1402, 12'sd1736}, {13'sd3109, 8'sd107, 12'sd1359}},
{{12'sd1237, 3'sd-2, 13'sd2727}, {13'sd-3678, 8'sd120, 10'sd-312}, {10'sd348, 8'sd-116, 12'sd1518}},
{{12'sd-1502, 10'sd459, 12'sd-2035}, {11'sd-799, 13'sd-2457, 11'sd-527}, {13'sd-2565, 12'sd-2028, 12'sd1310}},
{{14'sd4441, 11'sd880, 13'sd3777}, {12'sd1895, 10'sd308, 7'sd35}, {14'sd-4257, 14'sd-8133, 14'sd-4545}},
{{11'sd-530, 12'sd1042, 10'sd352}, {11'sd558, 13'sd2233, 13'sd3564}, {13'sd3293, 12'sd1476, 12'sd1389}},
{{12'sd1125, 12'sd-2011, 11'sd745}, {13'sd2084, 12'sd1190, 9'sd175}, {12'sd1909, 13'sd2241, 11'sd813}},
{{12'sd-1984, 13'sd2478, 13'sd3310}, {11'sd1006, 11'sd-1023, 8'sd79}, {14'sd4680, 12'sd1989, 13'sd2321}},
{{13'sd2874, 11'sd-536, 13'sd-2318}, {13'sd3201, 13'sd-2182, 12'sd-1948}, {12'sd-1128, 9'sd183, 10'sd-443}},
{{11'sd-854, 13'sd2121, 12'sd-1159}, {10'sd313, 8'sd-77, 12'sd1415}, {12'sd1217, 13'sd-2862, 10'sd-408}},
{{12'sd1928, 13'sd-3612, 13'sd-2466}, {11'sd-883, 11'sd874, 10'sd490}, {12'sd1733, 11'sd576, 11'sd932}},
{{14'sd-4470, 12'sd1349, 10'sd317}, {12'sd-1729, 13'sd-2548, 10'sd-324}, {12'sd1150, 13'sd-2056, 10'sd286}}},
{
{{11'sd-529, 12'sd2027, 10'sd470}, {12'sd-2015, 12'sd-1947, 13'sd-2540}, {13'sd-2585, 12'sd1028, 13'sd-2124}},
{{12'sd-1840, 12'sd-1170, 12'sd-1616}, {12'sd-1900, 12'sd-1123, 13'sd-2246}, {13'sd2174, 13'sd-2083, 13'sd-2153}},
{{12'sd-1882, 12'sd-1507, 13'sd-2998}, {12'sd1906, 12'sd-1796, 12'sd1550}, {12'sd-1537, 13'sd2440, 13'sd2077}},
{{13'sd2049, 11'sd-742, 12'sd1253}, {12'sd1589, 9'sd251, 12'sd-1962}, {12'sd-1608, 12'sd-1660, 10'sd-392}},
{{5'sd-15, 13'sd-2152, 12'sd-1788}, {12'sd1754, 12'sd1741, 12'sd1126}, {13'sd2252, 13'sd-2198, 12'sd1290}},
{{11'sd-712, 12'sd-1852, 13'sd-4008}, {13'sd-2226, 10'sd366, 12'sd-1080}, {11'sd598, 13'sd-2321, 13'sd-3617}},
{{13'sd2592, 13'sd-2683, 13'sd-2914}, {12'sd1702, 13'sd-2286, 14'sd-4863}, {12'sd1176, 12'sd1135, 14'sd-4596}},
{{13'sd-2296, 13'sd-2980, 11'sd-1007}, {12'sd-1847, 11'sd781, 12'sd1657}, {12'sd-2044, 13'sd-2860, 11'sd539}},
{{12'sd1869, 9'sd228, 13'sd2268}, {8'sd-73, 12'sd-1501, 13'sd2478}, {13'sd2083, 13'sd2416, 7'sd-58}},
{{13'sd2659, 12'sd-1473, 9'sd-235}, {12'sd1514, 9'sd-248, 13'sd2162}, {13'sd-2580, 13'sd-2138, 10'sd504}},
{{12'sd1472, 12'sd-1061, 12'sd1678}, {13'sd-2314, 13'sd2117, 12'sd-1455}, {13'sd-2392, 12'sd-2028, 12'sd1507}},
{{8'sd65, 8'sd-115, 12'sd1541}, {11'sd-689, 13'sd2588, 12'sd1581}, {6'sd-29, 12'sd1363, 12'sd-1805}},
{{13'sd2112, 13'sd3014, 10'sd-299}, {13'sd3083, 12'sd1762, 11'sd731}, {12'sd-1024, 13'sd-2914, 12'sd1592}},
{{12'sd-1601, 13'sd-2103, 11'sd940}, {11'sd908, 11'sd-654, 12'sd1723}, {10'sd-293, 12'sd-1538, 13'sd3094}},
{{12'sd-1525, 13'sd3876, 14'sd4825}, {10'sd494, 13'sd3378, 11'sd-560}, {13'sd-2265, 13'sd-2234, 13'sd-3378}},
{{10'sd490, 12'sd1180, 12'sd1840}, {13'sd3213, 9'sd250, 12'sd1386}, {11'sd854, 13'sd3779, 11'sd634}},
{{12'sd-1183, 8'sd-78, 13'sd2103}, {9'sd208, 12'sd1849, 12'sd1055}, {12'sd1814, 9'sd170, 11'sd564}},
{{10'sd-408, 11'sd-909, 9'sd146}, {12'sd1379, 13'sd-2170, 12'sd1724}, {13'sd3414, 12'sd-1815, 12'sd2013}},
{{12'sd-1399, 12'sd1461, 13'sd2809}, {12'sd1375, 12'sd1525, 12'sd1750}, {13'sd2475, 10'sd389, 11'sd-645}},
{{11'sd893, 12'sd1284, 10'sd271}, {12'sd-1154, 12'sd1893, 7'sd-56}, {13'sd-2128, 10'sd315, 11'sd983}},
{{11'sd550, 11'sd-920, 12'sd1700}, {10'sd-438, 11'sd-597, 12'sd-1045}, {10'sd-496, 12'sd1857, 12'sd-1663}},
{{13'sd2263, 13'sd-2355, 12'sd-1539}, {11'sd986, 3'sd-3, 13'sd2233}, {12'sd-1881, 12'sd-1455, 11'sd-992}},
{{11'sd-1002, 12'sd1420, 7'sd-54}, {13'sd-2388, 12'sd-1055, 12'sd-1985}, {12'sd-1192, 10'sd487, 11'sd-521}},
{{12'sd-1795, 12'sd-2032, 12'sd1294}, {11'sd590, 12'sd1026, 13'sd2909}, {13'sd2099, 12'sd-1287, 12'sd1685}},
{{11'sd761, 10'sd413, 11'sd825}, {13'sd-2111, 12'sd-1247, 11'sd-726}, {13'sd2943, 11'sd-842, 11'sd-563}},
{{13'sd2826, 10'sd-281, 13'sd2228}, {10'sd508, 13'sd2082, 12'sd1988}, {12'sd1892, 7'sd46, 13'sd-3020}},
{{9'sd-160, 11'sd689, 13'sd-3804}, {13'sd2697, 13'sd2407, 11'sd591}, {13'sd2431, 11'sd604, 13'sd-2211}},
{{13'sd2603, 10'sd468, 13'sd2480}, {10'sd-353, 13'sd-2254, 12'sd-1338}, {11'sd-683, 12'sd1103, 13'sd-2854}},
{{13'sd-2551, 11'sd716, 13'sd2495}, {11'sd-582, 12'sd1956, 12'sd1419}, {10'sd-450, 9'sd195, 11'sd957}},
{{9'sd251, 8'sd-123, 12'sd-1160}, {8'sd-125, 11'sd-600, 13'sd-2252}, {12'sd1037, 12'sd1341, 12'sd-1999}},
{{13'sd-2296, 13'sd-2956, 11'sd801}, {11'sd-699, 13'sd-2624, 12'sd-1341}, {12'sd-1919, 10'sd-404, 12'sd-1553}},
{{12'sd1499, 13'sd2417, 10'sd-502}, {12'sd-1803, 9'sd152, 13'sd2213}, {10'sd-375, 10'sd407, 13'sd-2597}},
{{13'sd-2258, 12'sd-1214, 10'sd288}, {13'sd-2166, 12'sd1675, 12'sd1863}, {12'sd1117, 13'sd-2743, 11'sd-996}},
{{13'sd-2197, 12'sd-1894, 11'sd-588}, {12'sd2047, 11'sd913, 10'sd-357}, {12'sd-1468, 12'sd1547, 12'sd1461}},
{{12'sd1104, 13'sd-3131, 13'sd2198}, {12'sd1404, 13'sd-2576, 12'sd1231}, {5'sd-12, 11'sd929, 13'sd3079}},
{{13'sd-2252, 12'sd-1027, 12'sd-1295}, {10'sd305, 13'sd-3023, 13'sd-2163}, {12'sd1810, 13'sd2084, 11'sd-604}},
{{12'sd1064, 13'sd-3212, 12'sd-1456}, {13'sd2136, 12'sd1635, 12'sd1427}, {11'sd-568, 9'sd-248, 13'sd-2130}},
{{12'sd1328, 13'sd-2591, 12'sd1658}, {12'sd1372, 12'sd-1453, 12'sd1500}, {13'sd2165, 10'sd-322, 13'sd3152}},
{{12'sd1516, 13'sd2205, 11'sd-811}, {12'sd1134, 13'sd-2413, 12'sd1560}, {13'sd-2547, 12'sd-1205, 12'sd1576}},
{{7'sd47, 6'sd-28, 12'sd-1249}, {13'sd-2507, 12'sd1975, 13'sd2088}, {11'sd868, 12'sd-1548, 11'sd-535}},
{{13'sd2739, 8'sd83, 12'sd-1544}, {12'sd-1721, 11'sd-657, 12'sd-1166}, {11'sd-773, 12'sd-1234, 12'sd-1362}},
{{13'sd-2487, 10'sd457, 12'sd1297}, {13'sd2255, 12'sd-1364, 9'sd132}, {12'sd1326, 13'sd-3015, 13'sd-3239}},
{{13'sd-2080, 13'sd2389, 13'sd-2501}, {12'sd-1602, 7'sd-45, 13'sd-2152}, {13'sd-3750, 13'sd-4046, 13'sd-3712}},
{{13'sd-2667, 11'sd-1016, 13'sd-3210}, {12'sd1551, 12'sd-1278, 9'sd-190}, {14'sd4762, 11'sd907, 14'sd-4629}},
{{13'sd2195, 11'sd-737, 11'sd-533}, {12'sd-1114, 12'sd-1634, 13'sd-2479}, {9'sd241, 12'sd1108, 13'sd2503}},
{{11'sd-848, 13'sd-3177, 13'sd-2311}, {12'sd-1977, 7'sd59, 13'sd2675}, {12'sd1600, 13'sd-2498, 13'sd2406}},
{{12'sd1809, 13'sd2200, 12'sd-1434}, {12'sd1790, 11'sd564, 12'sd-1395}, {12'sd2005, 12'sd-1817, 13'sd-2241}},
{{11'sd-565, 8'sd85, 12'sd1671}, {12'sd1670, 12'sd-1637, 12'sd1598}, {12'sd1475, 12'sd-1293, 13'sd2205}},
{{12'sd-2001, 12'sd1306, 10'sd489}, {10'sd411, 12'sd-1871, 13'sd-2113}, {12'sd1637, 11'sd685, 13'sd-4065}},
{{12'sd-1326, 9'sd164, 13'sd2284}, {9'sd-157, 10'sd459, 13'sd3765}, {13'sd2541, 12'sd1807, 11'sd689}},
{{11'sd989, 12'sd1259, 10'sd-315}, {13'sd-2342, 13'sd2509, 13'sd2400}, {7'sd63, 12'sd1791, 13'sd3827}},
{{12'sd-1362, 11'sd907, 12'sd-1314}, {13'sd-2281, 12'sd-1807, 12'sd-1500}, {13'sd-2245, 12'sd-1521, 11'sd908}},
{{11'sd983, 13'sd2290, 11'sd-971}, {11'sd903, 12'sd1988, 13'sd-2969}, {13'sd-2616, 12'sd-1437, 13'sd-3897}},
{{9'sd-181, 13'sd-2316, 12'sd-1409}, {12'sd-1304, 13'sd2084, 13'sd2083}, {11'sd555, 11'sd-842, 12'sd1728}},
{{13'sd2210, 12'sd1514, 13'sd-2549}, {13'sd2365, 11'sd-747, 12'sd1204}, {13'sd-2635, 11'sd944, 12'sd-1923}},
{{12'sd-1079, 12'sd-1700, 13'sd2324}, {11'sd753, 11'sd926, 12'sd-1040}, {13'sd-2780, 12'sd-1930, 13'sd-3044}},
{{12'sd1024, 14'sd4357, 13'sd3562}, {12'sd1364, 13'sd3439, 7'sd-34}, {14'sd-5099, 11'sd-936, 12'sd-2017}},
{{12'sd-1479, 13'sd2313, 12'sd1422}, {12'sd-1899, 12'sd1362, 13'sd3090}, {13'sd3504, 13'sd2702, 13'sd3738}},
{{13'sd2247, 12'sd-1658, 11'sd832}, {8'sd92, 11'sd-800, 11'sd974}, {12'sd-1963, 10'sd-501, 10'sd290}},
{{13'sd2090, 12'sd1090, 12'sd-1597}, {11'sd760, 10'sd-421, 12'sd1278}, {14'sd7543, 14'sd4997, 13'sd2171}},
{{13'sd2537, 13'sd2463, 12'sd1060}, {13'sd2387, 12'sd-2032, 13'sd2788}, {12'sd1277, 13'sd2374, 12'sd1121}},
{{12'sd1286, 11'sd706, 10'sd-322}, {12'sd-1073, 12'sd1407, 7'sd62}, {11'sd591, 11'sd-662, 12'sd-1878}},
{{13'sd-2656, 13'sd-2662, 13'sd-2427}, {9'sd-216, 12'sd-1832, 13'sd2171}, {10'sd-480, 12'sd-1234, 12'sd-1535}},
{{13'sd-2391, 13'sd-3429, 10'sd264}, {11'sd-873, 13'sd-2782, 11'sd596}, {10'sd325, 10'sd-400, 13'sd-2488}}},
{
{{13'sd-3065, 11'sd694, 13'sd-2344}, {12'sd-1598, 10'sd-422, 13'sd3254}, {12'sd1207, 13'sd-3138, 9'sd-245}},
{{12'sd-1844, 10'sd485, 12'sd-1416}, {11'sd904, 13'sd-2049, 12'sd1666}, {11'sd-856, 9'sd162, 12'sd-1369}},
{{12'sd-1024, 12'sd1705, 12'sd1583}, {13'sd-2245, 11'sd631, 13'sd2378}, {12'sd1024, 8'sd-65, 12'sd-1215}},
{{13'sd3326, 13'sd2819, 12'sd1519}, {11'sd-941, 9'sd214, 14'sd-4149}, {9'sd-190, 13'sd-2753, 12'sd-1570}},
{{13'sd2907, 14'sd5875, 14'sd6105}, {14'sd4524, 13'sd2858, 10'sd398}, {12'sd1720, 13'sd3756, 13'sd-2053}},
{{15'sd-10516, 11'sd-762, 12'sd-1576}, {14'sd-4126, 12'sd-1135, 12'sd1758}, {13'sd-2133, 13'sd-3592, 13'sd3856}},
{{12'sd-1598, 12'sd1470, 13'sd-2471}, {13'sd-3090, 14'sd-4472, 12'sd-1269}, {15'sd-11543, 15'sd-13506, 15'sd-9497}},
{{12'sd1680, 12'sd1303, 10'sd446}, {12'sd-1225, 10'sd-343, 12'sd-1201}, {13'sd-2682, 13'sd-3055, 13'sd-2117}},
{{13'sd-3065, 12'sd-1703, 10'sd370}, {12'sd-1396, 13'sd2713, 13'sd2669}, {13'sd-2892, 13'sd2511, 12'sd1240}},
{{12'sd1884, 13'sd2074, 12'sd1033}, {8'sd89, 12'sd-1338, 13'sd-2445}, {10'sd314, 13'sd-2901, 13'sd-3188}},
{{14'sd6523, 13'sd2914, 9'sd-153}, {12'sd1813, 10'sd-338, 13'sd-2679}, {13'sd-2455, 11'sd-637, 13'sd-2921}},
{{14'sd-5027, 12'sd1332, 13'sd3888}, {12'sd1258, 13'sd3437, 13'sd3930}, {14'sd4618, 13'sd3172, 13'sd3782}},
{{9'sd156, 12'sd-1211, 13'sd-3784}, {12'sd-1769, 13'sd-2378, 12'sd-1166}, {13'sd-2877, 14'sd-4529, 13'sd-3373}},
{{12'sd1379, 11'sd-607, 10'sd410}, {13'sd2951, 9'sd-243, 10'sd-495}, {12'sd1657, 12'sd1818, 13'sd-2084}},
{{14'sd6072, 14'sd6402, 15'sd14218}, {5'sd-10, 12'sd1549, 13'sd2361}, {11'sd713, 13'sd3039, 14'sd-4351}},
{{13'sd-3214, 13'sd-3943, 13'sd-2410}, {11'sd637, 12'sd1385, 10'sd-285}, {11'sd-942, 12'sd-1728, 13'sd2585}},
{{10'sd486, 13'sd-2113, 12'sd1394}, {10'sd410, 10'sd497, 12'sd-1082}, {13'sd2279, 13'sd3645, 11'sd-881}},
{{11'sd811, 8'sd121, 12'sd1351}, {12'sd-1321, 11'sd753, 13'sd-2957}, {12'sd-1069, 11'sd-711, 11'sd-628}},
{{10'sd-419, 8'sd-96, 11'sd847}, {11'sd1013, 13'sd-3779, 13'sd-2699}, {11'sd699, 12'sd-1734, 12'sd1465}},
{{12'sd-1201, 13'sd-2440, 11'sd-777}, {12'sd-1582, 11'sd-824, 10'sd429}, {12'sd1752, 11'sd555, 13'sd-2255}},
{{13'sd2712, 11'sd-946, 13'sd2750}, {11'sd-621, 12'sd-1600, 10'sd-421}, {10'sd307, 11'sd-544, 13'sd-2502}},
{{11'sd999, 13'sd2307, 12'sd-1245}, {12'sd-1538, 10'sd-358, 13'sd-4012}, {13'sd3096, 3'sd3, 12'sd-1420}},
{{10'sd-389, 12'sd1388, 12'sd1568}, {10'sd278, 13'sd2861, 13'sd2253}, {13'sd3387, 13'sd3897, 12'sd1749}},
{{13'sd-3061, 13'sd-3235, 13'sd-2145}, {12'sd1120, 13'sd2264, 10'sd-309}, {12'sd1076, 13'sd-2760, 12'sd-1306}},
{{14'sd4251, 11'sd808, 12'sd1190}, {13'sd2097, 10'sd312, 11'sd671}, {11'sd589, 13'sd-2382, 9'sd-191}},
{{12'sd1216, 13'sd3689, 11'sd931}, {12'sd-1490, 13'sd3363, 10'sd-487}, {12'sd2011, 11'sd-956, 13'sd2099}},
{{13'sd3431, 12'sd1204, 8'sd81}, {11'sd-512, 13'sd-3621, 13'sd-3085}, {13'sd-3928, 12'sd-1168, 11'sd-722}},
{{13'sd-3699, 11'sd-797, 12'sd1687}, {11'sd-807, 8'sd-67, 12'sd1981}, {11'sd-909, 11'sd837, 11'sd-925}},
{{14'sd4108, 13'sd3136, 14'sd4102}, {13'sd3035, 9'sd153, 12'sd-1475}, {13'sd3225, 13'sd-3574, 11'sd1018}},
{{11'sd-937, 12'sd-1965, 13'sd-2130}, {12'sd-1194, 11'sd967, 13'sd2355}, {12'sd-1230, 9'sd215, 11'sd-614}},
{{10'sd364, 6'sd-25, 12'sd-1917}, {11'sd-753, 12'sd-1568, 10'sd-337}, {13'sd3475, 9'sd224, 9'sd-159}},
{{12'sd-1240, 9'sd208, 13'sd3738}, {13'sd3098, 12'sd1122, 13'sd3199}, {12'sd-1198, 13'sd-2456, 13'sd2119}},
{{11'sd566, 13'sd-2434, 10'sd-340}, {11'sd-1012, 9'sd152, 13'sd-3052}, {13'sd-2086, 12'sd1516, 12'sd1653}},
{{12'sd-1518, 13'sd-2348, 11'sd821}, {9'sd-167, 13'sd2145, 11'sd738}, {12'sd-1764, 11'sd921, 11'sd910}},
{{13'sd-2976, 9'sd-150, 10'sd-418}, {13'sd-2335, 11'sd848, 13'sd-2506}, {13'sd3389, 13'sd2459, 13'sd3304}},
{{12'sd-2030, 11'sd-549, 9'sd209}, {10'sd506, 12'sd1674, 11'sd732}, {11'sd652, 11'sd533, 13'sd-3626}},
{{13'sd-3565, 13'sd-2896, 13'sd-2833}, {14'sd-4603, 10'sd-269, 12'sd1380}, {14'sd-5837, 12'sd1349, 10'sd417}},
{{12'sd1452, 13'sd3177, 10'sd-442}, {10'sd-398, 13'sd-2598, 13'sd-4078}, {14'sd-4823, 14'sd-6656, 14'sd-5749}},
{{13'sd2106, 12'sd2026, 9'sd-136}, {12'sd2003, 13'sd2232, 12'sd1950}, {13'sd-2238, 12'sd1025, 12'sd1359}},
{{12'sd1089, 9'sd168, 10'sd-292}, {12'sd-1605, 12'sd1745, 13'sd2474}, {12'sd-1138, 13'sd2346, 12'sd1213}},
{{10'sd-280, 13'sd-3131, 12'sd-1868}, {9'sd-245, 12'sd-1928, 14'sd-5313}, {13'sd-2373, 14'sd-4624, 14'sd-5722}},
{{14'sd4394, 13'sd3307, 10'sd420}, {13'sd2622, 13'sd2558, 12'sd1143}, {13'sd-2578, 13'sd-3940, 13'sd-3236}},
{{14'sd5410, 13'sd2104, 10'sd-331}, {13'sd2057, 11'sd-620, 14'sd-5698}, {14'sd-4715, 12'sd-1654, 11'sd-778}},
{{15'sd13659, 15'sd8263, 14'sd6761}, {14'sd8054, 12'sd1725, 12'sd1545}, {14'sd4150, 11'sd-963, 13'sd3270}},
{{13'sd-2825, 13'sd-2535, 12'sd-1404}, {13'sd-3391, 13'sd-2080, 13'sd2197}, {12'sd-1449, 13'sd-3063, 12'sd-1164}},
{{12'sd1458, 13'sd2817, 10'sd291}, {11'sd-917, 13'sd2808, 11'sd824}, {13'sd2124, 12'sd1137, 13'sd3585}},
{{14'sd-5305, 13'sd-2260, 14'sd-5127}, {11'sd-945, 13'sd-2492, 12'sd-1683}, {13'sd-3067, 11'sd-643, 10'sd305}},
{{13'sd3312, 13'sd2641, 10'sd271}, {12'sd-1574, 10'sd-446, 12'sd-1671}, {12'sd-1817, 11'sd-888, 13'sd-2498}},
{{14'sd-7218, 11'sd-513, 12'sd1067}, {14'sd-7200, 13'sd-3121, 10'sd-310}, {14'sd-6223, 12'sd-1156, 13'sd3895}},
{{14'sd-6445, 12'sd-1835, 13'sd-3737}, {13'sd-2727, 8'sd-67, 8'sd79}, {13'sd3324, 13'sd2212, 14'sd5183}},
{{13'sd2408, 12'sd-1202, 13'sd2262}, {13'sd2409, 11'sd-806, 13'sd-2230}, {14'sd5859, 12'sd2015, 12'sd1713}},
{{11'sd746, 12'sd-1697, 11'sd-864}, {9'sd135, 13'sd-2233, 13'sd2525}, {12'sd-1154, 10'sd-304, 11'sd755}},
{{13'sd3263, 13'sd2186, 12'sd1658}, {12'sd1367, 12'sd1787, 13'sd-2694}, {13'sd3338, 13'sd-2831, 12'sd-1778}},
{{11'sd913, 13'sd-2306, 13'sd-2722}, {11'sd-774, 11'sd532, 11'sd-1023}, {4'sd4, 9'sd254, 13'sd-3325}},
{{13'sd3458, 12'sd-1436, 13'sd-3301}, {11'sd762, 13'sd-2967, 13'sd-2985}, {14'sd-6021, 13'sd-4051, 15'sd-8622}},
{{13'sd-3685, 11'sd533, 13'sd-3603}, {11'sd988, 11'sd514, 11'sd-872}, {13'sd-2571, 12'sd1253, 11'sd599}},
{{15'sd11245, 13'sd3041, 11'sd657}, {13'sd2439, 12'sd-1532, 14'sd-5607}, {14'sd7128, 12'sd-1177, 14'sd-4292}},
{{12'sd-1857, 12'sd-1506, 10'sd398}, {12'sd1708, 11'sd-702, 12'sd-1331}, {13'sd3626, 10'sd-501, 13'sd-2496}},
{{12'sd-1349, 13'sd3284, 11'sd978}, {12'sd1348, 12'sd-1879, 12'sd1459}, {8'sd94, 12'sd-1680, 10'sd-449}},
{{14'sd-5537, 8'sd-69, 13'sd3542}, {13'sd-3792, 14'sd4120, 14'sd6999}, {14'sd-4747, 14'sd-5132, 12'sd-1437}},
{{10'sd-317, 13'sd2090, 8'sd114}, {13'sd-2777, 11'sd-747, 13'sd-3665}, {13'sd3490, 13'sd3512, 9'sd-190}},
{{13'sd-4051, 11'sd732, 12'sd1291}, {12'sd1369, 11'sd-944, 8'sd127}, {11'sd-773, 12'sd-1325, 13'sd-3392}},
{{11'sd871, 12'sd1256, 9'sd-255}, {8'sd-108, 13'sd-2437, 14'sd-4393}, {9'sd187, 8'sd-111, 13'sd-2515}},
{{11'sd587, 9'sd-190, 11'sd923}, {11'sd785, 13'sd2390, 13'sd2963}, {13'sd2156, 11'sd547, 10'sd432}}},
{
{{13'sd-2385, 9'sd240, 11'sd-991}, {11'sd961, 8'sd-93, 11'sd841}, {12'sd-1702, 11'sd966, 11'sd622}},
{{10'sd-452, 3'sd-2, 12'sd-1821}, {10'sd-306, 12'sd-1878, 12'sd1071}, {13'sd2357, 10'sd263, 11'sd965}},
{{12'sd-1984, 13'sd-2178, 5'sd9}, {13'sd2498, 11'sd-608, 11'sd822}, {13'sd-2221, 10'sd270, 12'sd2042}},
{{12'sd-1792, 13'sd-2152, 13'sd2322}, {12'sd1184, 12'sd1359, 13'sd-2064}, {12'sd-1880, 13'sd-2606, 12'sd-1566}},
{{13'sd3954, 9'sd188, 11'sd-676}, {13'sd3409, 13'sd2594, 13'sd2312}, {13'sd2100, 11'sd-813, 13'sd3226}},
{{9'sd207, 11'sd-797, 13'sd-3140}, {11'sd-850, 10'sd-329, 12'sd-1824}, {11'sd-729, 11'sd879, 12'sd1246}},
{{13'sd2719, 12'sd-1808, 12'sd1294}, {13'sd3001, 12'sd-1099, 12'sd-1440}, {12'sd-1910, 13'sd-3348, 13'sd-2125}},
{{12'sd1986, 11'sd-646, 12'sd-1651}, {12'sd-1094, 13'sd2254, 7'sd43}, {8'sd98, 10'sd465, 12'sd-1645}},
{{13'sd2416, 13'sd2246, 13'sd2391}, {11'sd621, 7'sd-56, 9'sd-238}, {12'sd-1535, 9'sd170, 12'sd1553}},
{{12'sd-1905, 11'sd740, 11'sd-940}, {12'sd-1744, 13'sd3074, 13'sd2233}, {13'sd-2702, 10'sd-308, 13'sd-2057}},
{{4'sd4, 13'sd-2116, 13'sd2230}, {12'sd-1640, 9'sd-168, 12'sd1866}, {12'sd-1083, 13'sd-2408, 12'sd-1427}},
{{13'sd2417, 11'sd605, 7'sd-50}, {10'sd274, 13'sd-2553, 12'sd1274}, {13'sd2072, 12'sd1744, 12'sd1698}},
{{13'sd2262, 13'sd2227, 10'sd-302}, {12'sd1151, 11'sd-896, 13'sd2240}, {12'sd1951, 13'sd-2397, 10'sd365}},
{{13'sd2474, 11'sd774, 12'sd-1554}, {12'sd-1971, 12'sd1051, 13'sd-2113}, {12'sd1593, 12'sd1594, 12'sd-1670}},
{{13'sd2707, 12'sd-1938, 13'sd3420}, {11'sd663, 12'sd1122, 12'sd1201}, {5'sd15, 11'sd690, 12'sd-1342}},
{{11'sd-1010, 13'sd2370, 12'sd1110}, {11'sd562, 12'sd1211, 10'sd261}, {12'sd1965, 12'sd-1790, 12'sd-1520}},
{{12'sd-1608, 13'sd-2113, 12'sd1654}, {12'sd1330, 13'sd2465, 12'sd1208}, {10'sd497, 12'sd-1628, 13'sd2497}},
{{12'sd1223, 13'sd3072, 13'sd3424}, {10'sd317, 10'sd-465, 12'sd-1313}, {10'sd-351, 10'sd411, 11'sd697}},
{{12'sd2014, 12'sd1043, 13'sd2421}, {7'sd37, 13'sd-2678, 12'sd1677}, {13'sd-2111, 11'sd564, 8'sd83}},
{{12'sd-1165, 12'sd1619, 12'sd1312}, {11'sd-949, 11'sd-524, 12'sd-1742}, {12'sd1489, 12'sd-1451, 12'sd1836}},
{{8'sd-87, 13'sd-2519, 13'sd-2422}, {12'sd1753, 12'sd-1094, 12'sd-1983}, {12'sd1928, 12'sd-1562, 12'sd1349}},
{{10'sd-326, 11'sd919, 12'sd-1933}, {9'sd-241, 7'sd-53, 12'sd1833}, {11'sd584, 10'sd-298, 11'sd-672}},
{{12'sd1645, 12'sd-1934, 12'sd1602}, {11'sd625, 12'sd-1482, 11'sd944}, {13'sd2161, 12'sd-1433, 12'sd-1645}},
{{13'sd-2126, 12'sd1966, 12'sd-1614}, {12'sd-1044, 12'sd-1755, 12'sd-1782}, {11'sd625, 10'sd414, 13'sd-2342}},
{{13'sd-2504, 13'sd2574, 12'sd-1630}, {11'sd632, 13'sd-2085, 13'sd2171}, {13'sd2260, 12'sd-1624, 12'sd-1615}},
{{12'sd2000, 12'sd1286, 10'sd-261}, {9'sd-250, 9'sd221, 12'sd-1851}, {12'sd1497, 10'sd-378, 12'sd1651}},
{{10'sd467, 12'sd-1399, 12'sd-1864}, {11'sd812, 13'sd-2280, 11'sd848}, {12'sd1903, 12'sd-1135, 12'sd1771}},
{{13'sd-2094, 11'sd958, 12'sd1655}, {12'sd-1348, 11'sd870, 13'sd2431}, {8'sd82, 9'sd-132, 12'sd-1132}},
{{10'sd269, 12'sd-1825, 10'sd-259}, {13'sd-2424, 13'sd-2899, 10'sd408}, {12'sd1997, 12'sd-1933, 13'sd2384}},
{{12'sd1876, 10'sd382, 12'sd-1922}, {11'sd-553, 12'sd-1453, 11'sd744}, {13'sd-2544, 12'sd1518, 6'sd-24}},
{{13'sd2774, 12'sd-1385, 11'sd-784}, {13'sd2495, 12'sd-2026, 12'sd1357}, {11'sd646, 9'sd157, 9'sd236}},
{{13'sd-2780, 13'sd2379, 10'sd-389}, {13'sd-2431, 12'sd1883, 13'sd2648}, {12'sd2034, 11'sd-1012, 11'sd-962}},
{{11'sd-743, 9'sd204, 12'sd1112}, {12'sd-1857, 7'sd63, 12'sd1924}, {13'sd2500, 12'sd-1487, 11'sd-1021}},
{{13'sd2403, 13'sd-2552, 13'sd2785}, {12'sd-1663, 11'sd-801, 12'sd-1812}, {9'sd-227, 12'sd-1465, 12'sd1752}},
{{13'sd2234, 13'sd-2891, 12'sd1370}, {13'sd-2331, 12'sd-1202, 9'sd-251}, {10'sd-323, 7'sd-41, 12'sd-1197}},
{{12'sd1419, 12'sd-1846, 8'sd98}, {10'sd368, 12'sd-1612, 12'sd-1883}, {11'sd895, 9'sd-171, 12'sd-1427}},
{{12'sd-1617, 13'sd-2827, 12'sd1139}, {11'sd-759, 9'sd158, 12'sd-1399}, {9'sd-199, 12'sd1079, 12'sd-1686}},
{{10'sd-451, 11'sd934, 12'sd1650}, {13'sd2292, 12'sd-1807, 12'sd1963}, {8'sd-92, 12'sd1690, 12'sd-1774}},
{{12'sd-1779, 10'sd460, 13'sd-2131}, {11'sd645, 13'sd-2636, 10'sd508}, {13'sd2620, 12'sd-1611, 12'sd1045}},
{{12'sd1242, 13'sd2680, 13'sd2093}, {7'sd-33, 11'sd959, 12'sd-1498}, {12'sd1996, 12'sd1292, 12'sd-1754}},
{{12'sd-1604, 13'sd2311, 10'sd502}, {13'sd3039, 11'sd553, 13'sd2194}, {13'sd2795, 11'sd917, 13'sd2812}},
{{9'sd222, 11'sd597, 10'sd-455}, {11'sd-803, 12'sd1376, 13'sd2131}, {13'sd2632, 11'sd655, 12'sd1341}},
{{9'sd-194, 11'sd633, 12'sd-1177}, {11'sd-768, 12'sd-1041, 12'sd-1312}, {12'sd-1623, 12'sd1295, 11'sd719}},
{{11'sd-747, 12'sd1684, 12'sd-1678}, {12'sd-1851, 12'sd-1871, 8'sd81}, {10'sd-376, 12'sd1214, 9'sd-131}},
{{10'sd-424, 9'sd-232, 12'sd-1758}, {11'sd1005, 12'sd1631, 12'sd1414}, {11'sd-625, 10'sd401, 8'sd-123}},
{{12'sd-1882, 12'sd1633, 13'sd-2076}, {11'sd885, 12'sd-1043, 13'sd2579}, {13'sd-2353, 12'sd1083, 12'sd1600}},
{{12'sd1560, 9'sd-216, 12'sd-1957}, {13'sd-2660, 12'sd1740, 8'sd97}, {12'sd1944, 13'sd-2872, 12'sd1888}},
{{10'sd-259, 11'sd-1018, 12'sd-1886}, {13'sd2643, 9'sd255, 11'sd1013}, {13'sd3011, 12'sd-1989, 12'sd-1305}},
{{13'sd-2530, 11'sd-779, 11'sd810}, {10'sd-377, 12'sd-1483, 12'sd-1447}, {13'sd-3092, 12'sd-1313, 11'sd548}},
{{7'sd-38, 11'sd-963, 12'sd-1832}, {12'sd-1668, 13'sd-3390, 9'sd-128}, {12'sd1452, 13'sd-2916, 12'sd1482}},
{{9'sd-252, 13'sd-2674, 13'sd2333}, {10'sd270, 12'sd2019, 13'sd2395}, {12'sd-1524, 10'sd-406, 12'sd-1103}},
{{11'sd-555, 12'sd2018, 12'sd-1950}, {9'sd-191, 10'sd497, 11'sd789}, {13'sd-2765, 13'sd-2296, 13'sd2297}},
{{11'sd890, 12'sd2038, 13'sd2142}, {10'sd474, 9'sd160, 12'sd-1144}, {12'sd1047, 10'sd272, 9'sd247}},
{{10'sd-402, 12'sd1459, 11'sd726}, {9'sd141, 12'sd1863, 12'sd1831}, {11'sd-562, 10'sd404, 13'sd2247}},
{{10'sd-481, 12'sd1960, 13'sd2938}, {9'sd-185, 11'sd-834, 12'sd-1285}, {13'sd-2100, 12'sd1880, 13'sd2090}},
{{12'sd-1792, 12'sd1799, 13'sd-3122}, {13'sd-2573, 8'sd113, 12'sd1589}, {12'sd1172, 12'sd1443, 10'sd309}},
{{13'sd2662, 9'sd171, 10'sd-286}, {12'sd1743, 12'sd1810, 12'sd1685}, {13'sd2393, 12'sd2016, 13'sd3228}},
{{12'sd-1269, 12'sd-1808, 10'sd-342}, {12'sd1035, 11'sd-612, 9'sd199}, {11'sd-594, 11'sd-709, 12'sd-1162}},
{{12'sd1677, 13'sd-2463, 13'sd2682}, {12'sd-1927, 12'sd1964, 13'sd-2264}, {10'sd483, 12'sd1400, 13'sd2614}},
{{11'sd988, 8'sd-118, 12'sd2036}, {13'sd2813, 13'sd-2615, 4'sd4}, {13'sd2499, 8'sd-88, 11'sd763}},
{{10'sd383, 10'sd382, 13'sd2251}, {12'sd1755, 11'sd566, 12'sd-1753}, {10'sd299, 13'sd2191, 12'sd-1767}},
{{11'sd-803, 12'sd-1509, 13'sd2383}, {13'sd-2150, 12'sd1179, 12'sd-1914}, {12'sd-1136, 12'sd-1537, 12'sd1168}},
{{13'sd2171, 13'sd-2902, 8'sd-67}, {8'sd64, 12'sd-1967, 12'sd-1689}, {12'sd-1215, 12'sd1094, 12'sd1653}},
{{13'sd-2479, 12'sd-1377, 12'sd-1981}, {3'sd3, 13'sd-2151, 10'sd-321}, {12'sd1276, 11'sd659, 11'sd783}}},
{
{{12'sd-1328, 10'sd273, 10'sd357}, {11'sd982, 11'sd-989, 13'sd2884}, {12'sd-1860, 12'sd-1630, 12'sd1756}},
{{12'sd-1526, 11'sd859, 11'sd-637}, {13'sd-2485, 11'sd-653, 10'sd-394}, {13'sd2258, 12'sd1074, 13'sd3040}},
{{6'sd-16, 12'sd-1422, 10'sd-374}, {10'sd303, 9'sd-130, 12'sd-1451}, {12'sd1769, 12'sd1205, 12'sd-1379}},
{{13'sd2950, 13'sd2903, 12'sd1241}, {13'sd2945, 13'sd-2048, 12'sd-1406}, {13'sd-2263, 11'sd714, 13'sd-2583}},
{{11'sd674, 12'sd1796, 12'sd1711}, {11'sd-886, 11'sd985, 13'sd2677}, {11'sd623, 12'sd1075, 10'sd427}},
{{11'sd570, 13'sd4042, 11'sd657}, {13'sd2728, 5'sd15, 11'sd-763}, {12'sd-1262, 9'sd207, 9'sd229}},
{{11'sd517, 12'sd2004, 12'sd1494}, {13'sd2796, 11'sd-762, 13'sd2087}, {12'sd1341, 13'sd-2787, 13'sd-3158}},
{{11'sd-776, 11'sd523, 11'sd712}, {11'sd-586, 11'sd-720, 12'sd-1945}, {13'sd-2266, 12'sd1208, 10'sd-352}},
{{12'sd1556, 13'sd-2154, 12'sd1218}, {13'sd-2775, 13'sd-2535, 8'sd-79}, {12'sd1264, 12'sd-1367, 12'sd1051}},
{{12'sd1973, 12'sd-1963, 11'sd-771}, {11'sd-595, 13'sd-2641, 13'sd-2364}, {12'sd-2038, 10'sd-327, 9'sd154}},
{{12'sd-1335, 12'sd-1822, 13'sd-2819}, {6'sd29, 11'sd899, 10'sd-488}, {13'sd-2935, 12'sd1195, 10'sd462}},
{{13'sd-2469, 10'sd445, 13'sd2826}, {12'sd1747, 12'sd-1047, 11'sd967}, {11'sd596, 12'sd1257, 11'sd-770}},
{{12'sd-1049, 11'sd690, 13'sd2141}, {13'sd2124, 12'sd1681, 13'sd2741}, {13'sd-2665, 13'sd2107, 13'sd3011}},
{{8'sd-73, 12'sd1735, 11'sd1007}, {12'sd1937, 11'sd-933, 12'sd1099}, {13'sd-2369, 12'sd1325, 12'sd1447}},
{{11'sd-853, 13'sd3047, 14'sd5848}, {12'sd1317, 12'sd-1301, 12'sd1468}, {11'sd-744, 12'sd1335, 11'sd-955}},
{{13'sd-2521, 13'sd2829, 11'sd907}, {12'sd-1849, 12'sd1907, 11'sd-882}, {9'sd212, 13'sd2205, 12'sd-1346}},
{{11'sd981, 12'sd-1952, 11'sd-618}, {12'sd1491, 12'sd-1465, 12'sd1310}, {11'sd1021, 8'sd91, 11'sd-550}},
{{12'sd-1254, 8'sd-113, 12'sd-1103}, {11'sd-756, 12'sd1593, 12'sd1620}, {10'sd-393, 12'sd1676, 12'sd1608}},
{{12'sd-1758, 11'sd-811, 12'sd-1464}, {12'sd1296, 12'sd1337, 10'sd-370}, {13'sd-2149, 13'sd2508, 12'sd-1669}},
{{13'sd2938, 13'sd-2163, 9'sd-185}, {11'sd944, 12'sd-1559, 12'sd-1214}, {13'sd3035, 11'sd-709, 12'sd1460}},
{{13'sd2376, 12'sd1534, 13'sd-2724}, {12'sd1247, 12'sd-1320, 13'sd-2531}, {13'sd-2434, 11'sd-732, 11'sd-861}},
{{11'sd991, 11'sd878, 11'sd964}, {11'sd712, 13'sd2359, 13'sd-2622}, {12'sd1254, 12'sd-1449, 12'sd1105}},
{{6'sd-19, 9'sd-220, 13'sd-2485}, {13'sd-2141, 13'sd2803, 9'sd223}, {12'sd1901, 10'sd-413, 12'sd1776}},
{{11'sd552, 12'sd1401, 12'sd1566}, {13'sd2501, 12'sd-1065, 12'sd-1483}, {10'sd336, 10'sd-326, 12'sd1777}},
{{12'sd-1807, 12'sd-1938, 12'sd1889}, {11'sd-776, 13'sd2589, 11'sd-539}, {10'sd491, 10'sd321, 12'sd-1610}},
{{13'sd2075, 12'sd-2039, 13'sd3139}, {12'sd1828, 12'sd1272, 8'sd-126}, {10'sd-307, 13'sd2706, 13'sd2234}},
{{12'sd-1440, 10'sd-416, 13'sd-3319}, {12'sd-1025, 8'sd-79, 12'sd1670}, {13'sd2155, 10'sd491, 12'sd-1885}},
{{13'sd-2218, 11'sd-1014, 13'sd3851}, {12'sd1445, 13'sd2080, 13'sd4004}, {12'sd-1816, 12'sd-1625, 12'sd-1401}},
{{9'sd-182, 13'sd-2622, 9'sd190}, {11'sd574, 12'sd-1420, 11'sd625}, {10'sd427, 11'sd968, 11'sd-890}},
{{12'sd-1027, 13'sd-2150, 12'sd-1215}, {11'sd818, 10'sd482, 9'sd-241}, {12'sd1044, 12'sd1026, 13'sd-2860}},
{{13'sd2871, 13'sd-2150, 10'sd-377}, {12'sd-1068, 11'sd849, 6'sd-31}, {12'sd-1561, 12'sd-1949, 12'sd-1801}},
{{12'sd1766, 12'sd1827, 11'sd-1010}, {11'sd657, 8'sd95, 12'sd1446}, {12'sd-1462, 13'sd-2422, 10'sd405}},
{{11'sd-725, 13'sd-2500, 7'sd55}, {11'sd600, 13'sd-2156, 12'sd-1776}, {12'sd-1932, 13'sd-2304, 12'sd1070}},
{{9'sd184, 9'sd172, 12'sd-1939}, {10'sd317, 12'sd-1117, 12'sd1257}, {13'sd2503, 13'sd2808, 12'sd1253}},
{{12'sd-1614, 12'sd-1664, 8'sd-119}, {12'sd1840, 13'sd2051, 11'sd-590}, {12'sd1181, 11'sd-578, 13'sd-2498}},
{{8'sd-67, 12'sd1385, 12'sd-1979}, {13'sd2911, 10'sd456, 12'sd-1329}, {12'sd1194, 7'sd-49, 11'sd986}},
{{12'sd1240, 13'sd2446, 11'sd-912}, {12'sd-1592, 13'sd2084, 12'sd-1061}, {13'sd4081, 11'sd-780, 12'sd1409}},
{{13'sd2149, 11'sd-531, 13'sd2512}, {11'sd772, 12'sd1108, 11'sd-758}, {13'sd3502, 12'sd1541, 10'sd-478}},
{{10'sd438, 12'sd-1882, 12'sd1674}, {13'sd2523, 13'sd-2243, 10'sd425}, {11'sd703, 11'sd639, 12'sd-1507}},
{{11'sd-988, 13'sd2667, 10'sd-376}, {10'sd-296, 10'sd-374, 13'sd2742}, {7'sd33, 11'sd-597, 13'sd2424}},
{{13'sd3395, 13'sd3038, 12'sd1302}, {13'sd3195, 13'sd-2312, 11'sd-720}, {10'sd505, 13'sd3336, 13'sd-2164}},
{{13'sd-2519, 13'sd-2230, 12'sd1492}, {10'sd412, 12'sd-1258, 11'sd729}, {13'sd-3032, 13'sd-3184, 12'sd-1687}},
{{10'sd-337, 13'sd-3475, 12'sd-1624}, {13'sd2825, 12'sd1343, 13'sd-2413}, {13'sd2273, 13'sd-2706, 12'sd-1037}},
{{11'sd-612, 13'sd-2099, 13'sd-2966}, {11'sd580, 13'sd2401, 12'sd1099}, {9'sd253, 13'sd-2353, 14'sd-4353}},
{{13'sd-2573, 12'sd1829, 12'sd1369}, {13'sd2371, 12'sd-1371, 13'sd2662}, {13'sd2553, 13'sd3276, 9'sd142}},
{{11'sd756, 13'sd2838, 11'sd649}, {11'sd-796, 13'sd2659, 13'sd-2094}, {9'sd-208, 11'sd760, 11'sd-535}},
{{13'sd3084, 12'sd1528, 9'sd162}, {12'sd1484, 13'sd2881, 12'sd-1986}, {12'sd1272, 12'sd1263, 12'sd1535}},
{{10'sd-486, 13'sd-3008, 9'sd-199}, {9'sd145, 13'sd2138, 12'sd1633}, {13'sd2503, 11'sd676, 12'sd-1647}},
{{12'sd-1208, 9'sd238, 13'sd2106}, {10'sd510, 10'sd-475, 12'sd-1431}, {12'sd-1426, 9'sd-128, 13'sd-2828}},
{{10'sd477, 13'sd3322, 9'sd236}, {11'sd-543, 12'sd-1234, 12'sd1755}, {10'sd361, 13'sd3236, 12'sd-1503}},
{{8'sd-90, 13'sd-2767, 11'sd-892}, {9'sd-139, 13'sd-2911, 12'sd1647}, {13'sd2241, 12'sd-1785, 12'sd-1118}},
{{12'sd-1826, 10'sd-437, 12'sd1990}, {12'sd-1662, 10'sd-386, 6'sd-27}, {12'sd-1723, 13'sd-3187, 13'sd-2914}},
{{12'sd-1497, 13'sd-2531, 12'sd-1264}, {13'sd-2061, 13'sd-2381, 11'sd927}, {14'sd-4268, 12'sd-1147, 13'sd-2371}},
{{12'sd1559, 12'sd1938, 11'sd-934}, {10'sd-368, 11'sd-563, 8'sd-127}, {11'sd865, 12'sd-1488, 13'sd-2399}},
{{12'sd1567, 13'sd2654, 12'sd1734}, {10'sd273, 10'sd-424, 13'sd3609}, {4'sd-7, 11'sd-606, 10'sd384}},
{{9'sd182, 9'sd154, 11'sd602}, {12'sd1286, 10'sd436, 11'sd999}, {12'sd1237, 12'sd1131, 11'sd837}},
{{13'sd2719, 11'sd-927, 12'sd1251}, {10'sd406, 12'sd-1166, 13'sd2813}, {14'sd-7111, 13'sd-3688, 12'sd1883}},
{{12'sd-1090, 12'sd1458, 13'sd2679}, {10'sd-485, 13'sd3307, 13'sd3764}, {8'sd127, 11'sd-657, 13'sd2196}},
{{13'sd-2137, 12'sd-1180, 13'sd2102}, {7'sd60, 7'sd-32, 12'sd1755}, {9'sd220, 13'sd2592, 11'sd644}},
{{13'sd2542, 9'sd133, 12'sd1701}, {12'sd-1080, 12'sd-1051, 13'sd3366}, {13'sd2674, 11'sd894, 13'sd3434}},
{{9'sd-129, 13'sd2981, 12'sd-1714}, {13'sd2677, 12'sd-1063, 13'sd2320}, {11'sd644, 12'sd1310, 13'sd2440}},
{{8'sd102, 13'sd2324, 12'sd-1473}, {11'sd-878, 12'sd-1794, 13'sd2322}, {12'sd1414, 10'sd-264, 10'sd-300}},
{{13'sd2971, 11'sd717, 11'sd-984}, {13'sd3367, 12'sd1064, 10'sd-301}, {11'sd661, 12'sd1652, 11'sd-997}},
{{10'sd-284, 13'sd-2392, 13'sd-3052}, {9'sd245, 9'sd-238, 11'sd-588}, {12'sd1284, 12'sd-1567, 11'sd-632}}},
{
{{12'sd1617, 11'sd551, 10'sd310}, {13'sd-2362, 12'sd1741, 11'sd912}, {12'sd1311, 12'sd-1458, 13'sd2203}},
{{13'sd-2739, 11'sd581, 9'sd252}, {13'sd-2479, 13'sd2555, 12'sd1824}, {8'sd101, 12'sd1080, 13'sd2795}},
{{12'sd-1063, 13'sd-2189, 12'sd1994}, {12'sd1611, 13'sd-2336, 12'sd1381}, {11'sd-719, 12'sd1237, 13'sd-2060}},
{{12'sd1933, 11'sd-684, 13'sd2285}, {13'sd2056, 12'sd1172, 12'sd1875}, {12'sd-1380, 13'sd2359, 13'sd2657}},
{{12'sd-1595, 13'sd-4073, 6'sd17}, {11'sd683, 13'sd-3867, 5'sd10}, {13'sd-2172, 12'sd-1398, 12'sd-2035}},
{{12'sd1048, 13'sd2596, 13'sd2720}, {12'sd-1337, 12'sd-1066, 12'sd1288}, {12'sd-1419, 12'sd-1539, 13'sd2774}},
{{12'sd-1878, 13'sd2299, 13'sd2557}, {11'sd-912, 10'sd432, 12'sd-1416}, {13'sd-3364, 12'sd1547, 12'sd-1719}},
{{8'sd86, 11'sd581, 13'sd-2081}, {9'sd-243, 11'sd771, 12'sd1212}, {13'sd-2323, 13'sd-2212, 12'sd1445}},
{{12'sd-1281, 13'sd-2665, 12'sd1229}, {7'sd-56, 11'sd-709, 11'sd662}, {11'sd825, 12'sd-1164, 12'sd-1761}},
{{13'sd2410, 12'sd1134, 13'sd-2405}, {11'sd-796, 9'sd168, 12'sd1439}, {13'sd-2207, 13'sd2418, 13'sd2354}},
{{12'sd-1929, 12'sd1530, 12'sd-1032}, {11'sd-633, 12'sd-1891, 13'sd-2801}, {13'sd2360, 10'sd427, 12'sd1118}},
{{13'sd-2988, 5'sd12, 13'sd2550}, {12'sd-1178, 12'sd1077, 11'sd-873}, {9'sd181, 9'sd213, 8'sd86}},
{{11'sd-867, 12'sd2038, 12'sd-1638}, {12'sd-1325, 10'sd401, 10'sd-382}, {11'sd660, 13'sd2474, 13'sd2398}},
{{13'sd2323, 12'sd1318, 12'sd-1619}, {12'sd1781, 10'sd350, 11'sd843}, {11'sd-860, 12'sd1445, 8'sd83}},
{{12'sd-1768, 11'sd-941, 13'sd2648}, {13'sd-2381, 12'sd1124, 11'sd-584}, {10'sd477, 11'sd863, 13'sd-3426}},
{{12'sd1229, 12'sd1156, 13'sd-3051}, {12'sd1538, 12'sd-1379, 9'sd-244}, {11'sd-783, 11'sd991, 13'sd-2093}},
{{12'sd1570, 12'sd-1855, 11'sd725}, {12'sd1588, 12'sd-1073, 11'sd-575}, {13'sd-2194, 13'sd2070, 11'sd733}},
{{12'sd-2009, 13'sd-2560, 11'sd587}, {11'sd887, 11'sd749, 12'sd1713}, {12'sd1056, 13'sd-2377, 10'sd-314}},
{{9'sd-223, 12'sd-1186, 8'sd105}, {12'sd1811, 13'sd-2394, 12'sd1320}, {12'sd2033, 9'sd223, 12'sd1318}},
{{12'sd-1362, 12'sd1613, 8'sd-113}, {10'sd328, 13'sd-2253, 13'sd-2172}, {9'sd236, 12'sd-1306, 13'sd-2451}},
{{12'sd-1174, 12'sd-1867, 12'sd-1071}, {12'sd1535, 13'sd-2255, 12'sd1374}, {12'sd1994, 13'sd-2803, 12'sd1472}},
{{13'sd2405, 13'sd-2299, 11'sd-707}, {13'sd2247, 11'sd-687, 12'sd1976}, {10'sd278, 12'sd1319, 12'sd-1485}},
{{13'sd2633, 13'sd-2401, 12'sd-1253}, {13'sd2251, 12'sd-1138, 12'sd-1857}, {12'sd1055, 11'sd-969, 13'sd2872}},
{{12'sd1384, 13'sd-2477, 13'sd-2442}, {12'sd1039, 13'sd2671, 9'sd232}, {12'sd-1807, 13'sd-2415, 12'sd1901}},
{{12'sd-1371, 11'sd550, 10'sd339}, {13'sd2789, 10'sd479, 12'sd1798}, {11'sd947, 13'sd-2401, 10'sd-426}},
{{12'sd-1524, 12'sd-1894, 10'sd-260}, {13'sd2443, 11'sd-994, 13'sd2457}, {13'sd2427, 10'sd-400, 13'sd2245}},
{{13'sd4033, 12'sd1156, 13'sd-2981}, {8'sd68, 13'sd-2589, 12'sd-1805}, {13'sd-3592, 6'sd26, 11'sd-777}},
{{11'sd939, 12'sd1101, 12'sd1550}, {12'sd-1268, 12'sd-1150, 13'sd2080}, {13'sd-2078, 10'sd-317, 13'sd-2646}},
{{13'sd2606, 12'sd1699, 10'sd485}, {12'sd1550, 11'sd-860, 11'sd-1009}, {11'sd-642, 11'sd855, 13'sd2060}},
{{12'sd1849, 12'sd1902, 13'sd-2448}, {12'sd-1951, 11'sd625, 8'sd-75}, {13'sd2437, 12'sd1594, 12'sd1693}},
{{9'sd224, 10'sd469, 11'sd932}, {12'sd-1431, 12'sd1301, 11'sd825}, {6'sd18, 10'sd-431, 11'sd-1013}},
{{12'sd-1194, 12'sd1993, 13'sd3223}, {8'sd64, 13'sd2464, 10'sd418}, {13'sd-2219, 13'sd3065, 13'sd2234}},
{{13'sd2359, 13'sd2766, 11'sd-829}, {13'sd-2599, 12'sd-1572, 8'sd-95}, {10'sd327, 12'sd1928, 11'sd739}},
{{13'sd-3379, 11'sd675, 12'sd-1416}, {11'sd-694, 13'sd2762, 12'sd-1341}, {10'sd340, 11'sd-705, 12'sd-1052}},
{{12'sd1058, 10'sd348, 9'sd196}, {10'sd-394, 7'sd41, 12'sd-1465}, {12'sd-1071, 12'sd1502, 11'sd-929}},
{{13'sd2817, 10'sd-277, 13'sd2114}, {12'sd-1331, 12'sd-1304, 13'sd-2472}, {13'sd2316, 12'sd1786, 11'sd543}},
{{12'sd1456, 14'sd4871, 13'sd3660}, {12'sd1416, 14'sd4295, 11'sd-789}, {12'sd-1497, 12'sd1144, 13'sd2215}},
{{13'sd-2520, 5'sd-9, 10'sd-353}, {12'sd2036, 5'sd-14, 12'sd1123}, {12'sd-1818, 13'sd2192, 11'sd619}},
{{12'sd1907, 11'sd-771, 12'sd1508}, {10'sd-423, 13'sd2477, 9'sd231}, {13'sd2592, 12'sd-1107, 12'sd1277}},
{{11'sd802, 10'sd488, 13'sd2183}, {13'sd2621, 13'sd-2211, 11'sd773}, {11'sd601, 12'sd1027, 12'sd-1338}},
{{12'sd-1910, 12'sd-1226, 13'sd-2521}, {12'sd-1419, 13'sd-2892, 9'sd-136}, {12'sd-1153, 12'sd1932, 11'sd902}},
{{10'sd-286, 13'sd-2171, 11'sd893}, {11'sd941, 13'sd-2233, 12'sd-1558}, {11'sd-732, 12'sd-1370, 13'sd2550}},
{{10'sd357, 13'sd2270, 12'sd-1389}, {12'sd1352, 12'sd1715, 13'sd-3451}, {10'sd-492, 9'sd-157, 13'sd-3528}},
{{14'sd5518, 12'sd1388, 12'sd1762}, {13'sd3123, 12'sd1571, 13'sd2674}, {11'sd-513, 12'sd1797, 10'sd-336}},
{{13'sd-2676, 12'sd-1048, 12'sd1501}, {8'sd123, 7'sd-51, 9'sd180}, {12'sd-1305, 12'sd1641, 12'sd-1906}},
{{11'sd-720, 12'sd1351, 10'sd465}, {12'sd-1405, 12'sd-1231, 13'sd2696}, {10'sd-399, 12'sd-1745, 11'sd-877}},
{{12'sd1692, 13'sd2062, 13'sd2355}, {6'sd-21, 12'sd2014, 12'sd1299}, {13'sd-2752, 13'sd2060, 10'sd-318}},
{{7'sd42, 11'sd-869, 12'sd1199}, {12'sd-1053, 13'sd-2223, 12'sd-1939}, {12'sd1474, 11'sd991, 9'sd-222}},
{{11'sd-727, 13'sd2908, 12'sd2028}, {7'sd56, 12'sd1477, 12'sd-1727}, {9'sd232, 12'sd-1485, 12'sd-1375}},
{{13'sd2327, 13'sd3908, 13'sd-2434}, {13'sd2290, 13'sd2451, 10'sd-433}, {11'sd-850, 12'sd-1104, 11'sd648}},
{{11'sd-773, 13'sd-2117, 13'sd-3281}, {13'sd-2578, 13'sd2330, 3'sd2}, {11'sd841, 10'sd-434, 10'sd292}},
{{12'sd1426, 13'sd-2083, 8'sd-127}, {12'sd1513, 13'sd-2477, 12'sd-1452}, {12'sd1148, 12'sd1606, 12'sd1076}},
{{10'sd466, 13'sd2411, 11'sd905}, {11'sd-624, 11'sd-530, 12'sd1919}, {13'sd3253, 12'sd1466, 12'sd-1892}},
{{10'sd432, 13'sd2294, 11'sd-693}, {11'sd560, 11'sd714, 10'sd-432}, {12'sd1114, 13'sd-2746, 11'sd627}},
{{12'sd1593, 10'sd-299, 11'sd764}, {11'sd642, 9'sd205, 11'sd-995}, {12'sd1156, 12'sd1273, 13'sd-2311}},
{{12'sd1299, 13'sd2371, 12'sd1426}, {11'sd912, 12'sd1828, 11'sd919}, {11'sd564, 11'sd1007, 10'sd-454}},
{{14'sd5183, 10'sd-267, 13'sd-3136}, {12'sd-1985, 12'sd1350, 13'sd-2414}, {13'sd2888, 7'sd-48, 13'sd-2320}},
{{14'sd-4362, 12'sd-1919, 12'sd1089}, {11'sd-924, 11'sd-732, 13'sd-2681}, {10'sd315, 11'sd-1010, 12'sd-1082}},
{{12'sd-1796, 12'sd1524, 11'sd719}, {12'sd-1811, 12'sd-1420, 12'sd1507}, {11'sd-910, 12'sd1370, 12'sd1830}},
{{13'sd-2541, 10'sd446, 13'sd2575}, {12'sd-1299, 12'sd-1247, 12'sd-1618}, {12'sd-1055, 12'sd1061, 7'sd47}},
{{12'sd-1193, 12'sd1862, 12'sd-1237}, {11'sd-581, 13'sd-2456, 10'sd-264}, {9'sd-228, 13'sd2143, 11'sd760}},
{{13'sd-2387, 8'sd-112, 13'sd2367}, {11'sd-932, 12'sd1790, 12'sd-1813}, {12'sd1231, 12'sd1755, 8'sd68}},
{{9'sd252, 7'sd53, 11'sd588}, {11'sd943, 10'sd-379, 12'sd-1028}, {12'sd-1687, 10'sd393, 13'sd2516}},
{{11'sd-1023, 12'sd1065, 10'sd468}, {11'sd-604, 9'sd139, 12'sd-1792}, {12'sd-1844, 9'sd-237, 13'sd2225}}},
{
{{13'sd2964, 12'sd1469, 11'sd-660}, {8'sd-84, 12'sd-1302, 13'sd2058}, {13'sd2762, 12'sd1075, 12'sd-1565}},
{{13'sd2345, 10'sd335, 11'sd-789}, {11'sd-1006, 11'sd-542, 13'sd3044}, {12'sd1134, 9'sd-151, 12'sd-1349}},
{{8'sd103, 10'sd269, 11'sd-768}, {12'sd1119, 11'sd-871, 13'sd-2699}, {12'sd1326, 13'sd-2130, 12'sd-1504}},
{{11'sd-690, 6'sd19, 10'sd442}, {12'sd1532, 8'sd116, 9'sd-232}, {13'sd-2130, 12'sd1067, 11'sd696}},
{{13'sd-3794, 14'sd-4912, 10'sd-324}, {13'sd-2756, 14'sd-4152, 13'sd-3908}, {11'sd-985, 13'sd-2562, 13'sd-2647}},
{{11'sd902, 13'sd2397, 12'sd1299}, {12'sd1211, 13'sd-2261, 11'sd855}, {12'sd-1986, 12'sd-1833, 11'sd-734}},
{{13'sd-2977, 12'sd-2047, 10'sd318}, {12'sd-1350, 12'sd1910, 13'sd2138}, {11'sd874, 13'sd2768, 12'sd1428}},
{{13'sd2220, 11'sd526, 11'sd949}, {11'sd721, 12'sd1604, 10'sd-288}, {12'sd-1788, 13'sd-2050, 13'sd-2158}},
{{12'sd-1652, 12'sd-1339, 13'sd2214}, {13'sd2058, 9'sd206, 13'sd2483}, {11'sd-655, 12'sd-1635, 11'sd-929}},
{{8'sd104, 13'sd2632, 12'sd-1133}, {13'sd-2387, 9'sd-140, 11'sd-536}, {13'sd-2792, 8'sd-69, 12'sd1588}},
{{12'sd1424, 12'sd1304, 11'sd-971}, {12'sd1598, 13'sd2138, 10'sd455}, {11'sd-982, 13'sd2757, 13'sd-2633}},
{{12'sd1152, 11'sd801, 9'sd-228}, {12'sd-2015, 11'sd694, 9'sd-231}, {11'sd-756, 13'sd-2422, 11'sd-679}},
{{11'sd876, 10'sd421, 11'sd720}, {11'sd-830, 12'sd1437, 12'sd1950}, {13'sd2724, 11'sd679, 13'sd2453}},
{{10'sd263, 12'sd-1154, 12'sd-1947}, {9'sd-167, 12'sd-1688, 10'sd498}, {11'sd724, 9'sd170, 11'sd892}},
{{15'sd-8451, 14'sd-4806, 13'sd-2206}, {15'sd-10108, 14'sd-5812, 14'sd-6008}, {14'sd-6413, 14'sd-5434, 10'sd-324}},
{{11'sd861, 12'sd1547, 4'sd5}, {12'sd1835, 13'sd2386, 10'sd-478}, {14'sd4606, 13'sd3292, 13'sd2085}},
{{12'sd1995, 12'sd1998, 11'sd942}, {13'sd-2238, 11'sd516, 10'sd-345}, {12'sd-1129, 11'sd933, 12'sd-1386}},
{{12'sd1231, 12'sd-1307, 11'sd-665}, {13'sd-2406, 13'sd-2454, 12'sd-1099}, {10'sd271, 12'sd2046, 12'sd-1143}},
{{12'sd1567, 13'sd-2399, 10'sd-449}, {12'sd1407, 11'sd702, 13'sd2488}, {13'sd-2790, 11'sd-660, 12'sd-1337}},
{{13'sd-2933, 9'sd155, 11'sd-923}, {11'sd-809, 13'sd-2648, 13'sd2435}, {12'sd-1439, 12'sd1633, 12'sd1231}},
{{13'sd-3090, 10'sd-306, 11'sd1015}, {13'sd-2988, 12'sd1636, 13'sd-2197}, {8'sd-81, 10'sd-305, 12'sd1583}},
{{12'sd-1227, 12'sd1355, 8'sd94}, {11'sd-1006, 11'sd-915, 11'sd-841}, {12'sd1811, 12'sd1074, 11'sd903}},
{{11'sd521, 13'sd2643, 12'sd1147}, {12'sd-1599, 11'sd-778, 11'sd807}, {10'sd451, 13'sd-2434, 12'sd1807}},
{{12'sd-1074, 12'sd-1457, 12'sd-1891}, {13'sd2175, 13'sd2198, 11'sd849}, {11'sd-978, 11'sd-716, 12'sd1360}},
{{11'sd621, 13'sd2972, 12'sd1728}, {13'sd2812, 12'sd1086, 12'sd1055}, {11'sd861, 13'sd2447, 11'sd760}},
{{11'sd-725, 12'sd1950, 12'sd1781}, {3'sd2, 13'sd2505, 13'sd2483}, {12'sd1126, 12'sd-2020, 12'sd-1793}},
{{14'sd7349, 14'sd4582, 13'sd2968}, {15'sd9020, 14'sd4610, 12'sd1266}, {14'sd6614, 12'sd1438, 11'sd-801}},
{{10'sd-422, 13'sd-3387, 10'sd-488}, {13'sd-3366, 13'sd-2240, 10'sd454}, {13'sd-3768, 10'sd-381, 13'sd-2800}},
{{13'sd2748, 12'sd-1891, 9'sd158}, {11'sd-630, 9'sd227, 8'sd124}, {12'sd1106, 11'sd688, 12'sd-1642}},
{{12'sd-1398, 12'sd1792, 12'sd-2025}, {12'sd1592, 8'sd68, 12'sd1293}, {13'sd2640, 9'sd-225, 13'sd-2502}},
{{11'sd-688, 13'sd-2547, 11'sd951}, {11'sd-691, 13'sd-2102, 12'sd1440}, {12'sd-1359, 10'sd502, 12'sd1213}},
{{12'sd1105, 11'sd928, 13'sd3336}, {11'sd879, 10'sd-472, 12'sd-1730}, {13'sd2598, 11'sd605, 11'sd-838}},
{{11'sd919, 12'sd-1748, 13'sd2783}, {10'sd386, 11'sd-984, 12'sd1669}, {12'sd-1440, 13'sd2067, 13'sd-2127}},
{{9'sd239, 13'sd-2813, 13'sd-3443}, {11'sd-883, 13'sd2857, 12'sd1754}, {13'sd-2180, 13'sd2400, 12'sd1441}},
{{13'sd-2554, 12'sd1691, 12'sd-1767}, {12'sd-1837, 13'sd-2051, 9'sd-162}, {12'sd-1439, 11'sd581, 13'sd3043}},
{{11'sd594, 12'sd1982, 10'sd-284}, {9'sd-221, 13'sd-2700, 13'sd2139}, {10'sd-293, 13'sd-2546, 12'sd1660}},
{{10'sd401, 9'sd-239, 11'sd907}, {13'sd3534, 13'sd2896, 11'sd650}, {12'sd1302, 13'sd2831, 12'sd1512}},
{{12'sd2008, 12'sd1909, 12'sd-1380}, {11'sd928, 12'sd1046, 13'sd2463}, {11'sd592, 8'sd119, 11'sd-609}},
{{12'sd-1360, 12'sd1802, 11'sd-990}, {12'sd-1059, 11'sd-877, 11'sd978}, {8'sd112, 13'sd2055, 9'sd166}},
{{10'sd-313, 9'sd192, 13'sd-2651}, {12'sd-1860, 11'sd-795, 13'sd-2197}, {12'sd-1774, 8'sd91, 12'sd1695}},
{{10'sd-451, 9'sd220, 8'sd118}, {12'sd-1878, 10'sd-439, 10'sd257}, {11'sd-513, 10'sd-426, 12'sd1043}},
{{13'sd2750, 10'sd-417, 13'sd-2467}, {12'sd-1965, 13'sd2195, 11'sd988}, {8'sd108, 13'sd2683, 12'sd1952}},
{{11'sd996, 13'sd3874, 12'sd1592}, {11'sd-921, 12'sd2047, 9'sd-163}, {11'sd-961, 12'sd1241, 9'sd-243}},
{{14'sd5494, 13'sd4031, 14'sd4204}, {14'sd5850, 13'sd2770, 12'sd1269}, {14'sd8050, 14'sd7747, 12'sd1969}},
{{11'sd-876, 12'sd-1867, 11'sd514}, {12'sd1860, 11'sd600, 12'sd1417}, {13'sd2743, 13'sd2510, 13'sd2193}},
{{13'sd-2696, 12'sd-1532, 11'sd794}, {11'sd809, 11'sd872, 7'sd49}, {12'sd1763, 11'sd801, 11'sd-658}},
{{13'sd3514, 10'sd456, 12'sd-1838}, {13'sd3387, 12'sd1910, 12'sd1628}, {10'sd-415, 10'sd312, 12'sd-2021}},
{{9'sd142, 13'sd-2283, 11'sd-810}, {12'sd-1545, 11'sd728, 13'sd-3216}, {11'sd533, 12'sd-1311, 12'sd2025}},
{{12'sd1763, 13'sd-2359, 10'sd-256}, {10'sd-299, 6'sd16, 13'sd-2717}, {10'sd263, 12'sd1588, 12'sd-1623}},
{{12'sd-2028, 13'sd-2079, 13'sd2896}, {13'sd-2502, 13'sd-2666, 13'sd-2334}, {12'sd-1099, 13'sd-2871, 12'sd-1564}},
{{13'sd-3123, 12'sd-1155, 12'sd1236}, {13'sd-3873, 12'sd1755, 12'sd1241}, {13'sd-2496, 11'sd826, 12'sd-1759}},
{{12'sd1291, 8'sd65, 13'sd-2393}, {11'sd-531, 12'sd1123, 13'sd-2261}, {11'sd-626, 12'sd1692, 9'sd-229}},
{{13'sd-2942, 12'sd-1872, 11'sd-929}, {10'sd-495, 11'sd-731, 11'sd-773}, {12'sd-1973, 12'sd-1200, 11'sd-792}},
{{12'sd-1672, 13'sd2553, 12'sd1131}, {12'sd-1611, 10'sd-270, 11'sd-739}, {13'sd2284, 13'sd2467, 12'sd1541}},
{{11'sd871, 10'sd-501, 13'sd-2350}, {11'sd965, 12'sd-1238, 10'sd372}, {13'sd-2907, 10'sd306, 10'sd305}},
{{12'sd1301, 11'sd-954, 12'sd1067}, {13'sd-2664, 8'sd100, 12'sd-1547}, {13'sd-2227, 12'sd-1936, 13'sd2735}},
{{11'sd-888, 13'sd-2813, 13'sd2868}, {13'sd-3607, 12'sd1547, 12'sd1929}, {14'sd-4165, 12'sd1569, 13'sd2275}},
{{13'sd-2881, 10'sd-375, 12'sd-1990}, {11'sd-612, 12'sd1602, 12'sd-1238}, {10'sd461, 13'sd-2688, 13'sd-2657}},
{{13'sd2252, 12'sd-1697, 12'sd-1785}, {11'sd951, 13'sd-2198, 12'sd-1643}, {13'sd-2445, 11'sd591, 12'sd-1866}},
{{12'sd-1879, 12'sd-1159, 13'sd-3380}, {12'sd1988, 13'sd2099, 9'sd186}, {13'sd-2561, 12'sd-1827, 11'sd666}},
{{9'sd199, 9'sd233, 13'sd2257}, {12'sd-1064, 12'sd1183, 12'sd1704}, {13'sd-2693, 10'sd-336, 13'sd-2481}},
{{11'sd-525, 11'sd968, 8'sd125}, {13'sd-2515, 12'sd-1502, 11'sd883}, {11'sd-677, 12'sd-1326, 10'sd298}},
{{1'sd0, 12'sd1356, 12'sd1135}, {13'sd-2823, 12'sd1795, 13'sd2063}, {9'sd228, 12'sd-1253, 11'sd-824}},
{{11'sd-718, 13'sd-2340, 11'sd-662}, {11'sd914, 12'sd1973, 13'sd-2864}, {13'sd-2134, 8'sd88, 9'sd-218}}},
{
{{13'sd2450, 13'sd-2473, 13'sd2388}, {12'sd-1118, 13'sd2059, 12'sd-1871}, {11'sd-895, 12'sd-1979, 11'sd818}},
{{12'sd-1656, 13'sd2118, 13'sd-2070}, {9'sd130, 12'sd-1429, 12'sd-1517}, {11'sd-923, 9'sd227, 12'sd1559}},
{{11'sd717, 12'sd1280, 11'sd-517}, {10'sd434, 6'sd-19, 12'sd-1607}, {12'sd1499, 12'sd1315, 13'sd-2348}},
{{12'sd1499, 12'sd-1922, 11'sd617}, {13'sd-2841, 12'sd-1756, 13'sd2315}, {10'sd483, 13'sd-2865, 10'sd-320}},
{{13'sd-3249, 12'sd-1949, 13'sd-2620}, {13'sd-2735, 13'sd-3326, 7'sd-36}, {11'sd-731, 13'sd-2540, 8'sd90}},
{{10'sd289, 13'sd2378, 13'sd2636}, {7'sd50, 12'sd-1404, 12'sd1257}, {13'sd2162, 12'sd1413, 12'sd-1648}},
{{12'sd-1576, 13'sd-2149, 13'sd2337}, {12'sd-1396, 12'sd1444, 8'sd116}, {12'sd-1113, 12'sd1510, 11'sd550}},
{{13'sd2424, 13'sd2271, 12'sd-1283}, {12'sd-1452, 12'sd-1387, 10'sd-370}, {13'sd-2587, 11'sd-691, 12'sd1185}},
{{13'sd-2960, 6'sd-31, 13'sd-2431}, {13'sd2514, 11'sd736, 12'sd-1506}, {13'sd-2589, 9'sd131, 6'sd19}},
{{11'sd878, 13'sd2056, 11'sd-781}, {12'sd-1927, 10'sd-375, 10'sd-467}, {13'sd2435, 12'sd-1051, 11'sd901}},
{{13'sd2073, 12'sd-1858, 10'sd-355}, {10'sd349, 10'sd459, 10'sd-506}, {12'sd1365, 13'sd-2711, 12'sd1531}},
{{12'sd-1837, 10'sd279, 11'sd-617}, {11'sd-553, 11'sd-638, 12'sd-1695}, {12'sd-1593, 10'sd-476, 12'sd1515}},
{{10'sd-309, 12'sd1316, 12'sd1421}, {12'sd1599, 12'sd1756, 8'sd-94}, {11'sd924, 11'sd808, 11'sd687}},
{{10'sd390, 8'sd105, 12'sd1494}, {12'sd-1450, 12'sd-1973, 12'sd1594}, {11'sd904, 12'sd-1276, 12'sd-2047}},
{{11'sd969, 9'sd185, 10'sd-490}, {11'sd-578, 13'sd-2969, 13'sd-2471}, {14'sd-4421, 13'sd-2981, 7'sd-44}},
{{10'sd-510, 12'sd1252, 12'sd1901}, {12'sd1926, 12'sd-1135, 12'sd1319}, {12'sd-1518, 13'sd2056, 12'sd-1683}},
{{11'sd-648, 13'sd2208, 8'sd-77}, {11'sd-793, 12'sd1064, 12'sd1448}, {13'sd2929, 12'sd-1900, 12'sd1698}},
{{13'sd-3427, 12'sd1142, 8'sd-92}, {12'sd-1908, 12'sd-1278, 10'sd-381}, {13'sd-3820, 10'sd-287, 11'sd783}},
{{13'sd-2287, 10'sd484, 13'sd-2302}, {11'sd-903, 12'sd1881, 12'sd1643}, {11'sd894, 11'sd605, 12'sd1570}},
{{13'sd2810, 13'sd2974, 13'sd2058}, {13'sd2184, 13'sd-2300, 13'sd2679}, {13'sd2178, 13'sd-2388, 11'sd608}},
{{12'sd2037, 12'sd1888, 11'sd680}, {11'sd825, 12'sd1777, 13'sd-2247}, {13'sd-2386, 13'sd-2564, 11'sd897}},
{{4'sd6, 12'sd1092, 12'sd1803}, {12'sd1135, 12'sd-1879, 13'sd2308}, {12'sd-1328, 10'sd-508, 11'sd936}},
{{9'sd-134, 13'sd-2281, 13'sd2102}, {8'sd104, 10'sd-403, 11'sd883}, {12'sd1863, 12'sd-1311, 12'sd1193}},
{{12'sd1206, 12'sd1114, 9'sd-198}, {10'sd-315, 9'sd134, 13'sd2059}, {9'sd-155, 12'sd-1090, 12'sd1486}},
{{12'sd-1031, 10'sd273, 12'sd-1612}, {12'sd-1781, 12'sd-1157, 11'sd863}, {13'sd2345, 7'sd63, 10'sd-506}},
{{12'sd1030, 11'sd717, 12'sd1253}, {13'sd-2097, 12'sd-1097, 13'sd-2961}, {11'sd621, 9'sd-163, 12'sd-1379}},
{{12'sd-1262, 13'sd-2221, 13'sd2175}, {13'sd-2769, 11'sd-700, 12'sd-1244}, {12'sd-2030, 13'sd-2321, 12'sd-1596}},
{{8'sd127, 13'sd-2408, 11'sd914}, {10'sd465, 12'sd-1530, 12'sd1508}, {13'sd-2811, 12'sd1556, 12'sd-1429}},
{{13'sd2823, 12'sd-1989, 12'sd-1816}, {13'sd-2442, 13'sd2421, 12'sd-1206}, {13'sd-2250, 13'sd-2097, 10'sd-323}},
{{7'sd35, 10'sd397, 12'sd1291}, {12'sd1833, 9'sd-141, 12'sd1241}, {13'sd-2420, 10'sd279, 11'sd686}},
{{12'sd1717, 11'sd-845, 12'sd-1904}, {12'sd1668, 12'sd1139, 10'sd-421}, {13'sd2162, 13'sd2675, 13'sd2088}},
{{11'sd987, 13'sd2796, 12'sd-1114}, {11'sd-859, 10'sd290, 12'sd-1895}, {11'sd736, 9'sd-140, 10'sd292}},
{{11'sd661, 13'sd2289, 13'sd-2203}, {12'sd-1453, 11'sd686, 9'sd164}, {11'sd-812, 13'sd2109, 11'sd-1015}},
{{11'sd-777, 12'sd1352, 11'sd-689}, {13'sd-2138, 11'sd817, 13'sd-2239}, {11'sd-826, 7'sd42, 11'sd681}},
{{13'sd2564, 13'sd2889, 12'sd2021}, {12'sd-2006, 12'sd-1691, 12'sd-1473}, {13'sd2877, 12'sd-1058, 11'sd-708}},
{{9'sd-181, 13'sd-2214, 11'sd-548}, {9'sd153, 12'sd-1683, 13'sd2319}, {11'sd-830, 11'sd-698, 12'sd-1703}},
{{11'sd-565, 14'sd4098, 13'sd2933}, {11'sd-667, 12'sd1121, 13'sd3404}, {13'sd3685, 12'sd1484, 13'sd2804}},
{{11'sd-750, 13'sd-3019, 10'sd-466}, {12'sd-1458, 10'sd303, 11'sd633}, {9'sd157, 12'sd2040, 12'sd-1427}},
{{13'sd2316, 11'sd789, 12'sd1791}, {10'sd404, 10'sd-401, 12'sd-1384}, {5'sd10, 9'sd214, 10'sd-483}},
{{11'sd-772, 12'sd1217, 12'sd-1518}, {10'sd269, 13'sd-2430, 12'sd1124}, {5'sd-12, 13'sd-2196, 7'sd-51}},
{{11'sd978, 11'sd-723, 12'sd1306}, {8'sd-120, 13'sd2056, 10'sd263}, {11'sd-790, 7'sd-34, 12'sd-1411}},
{{12'sd1488, 8'sd-78, 11'sd999}, {13'sd-3117, 13'sd-2560, 11'sd684}, {11'sd-961, 9'sd-255, 13'sd-2129}},
{{12'sd1561, 12'sd1894, 12'sd1348}, {9'sd-239, 11'sd643, 9'sd-197}, {13'sd-2144, 12'sd-1354, 12'sd1491}},
{{11'sd876, 12'sd-1765, 13'sd3800}, {12'sd-1260, 8'sd109, 13'sd2375}, {12'sd1561, 11'sd-872, 12'sd-1812}},
{{12'sd1149, 10'sd-477, 10'sd486}, {12'sd1284, 7'sd62, 13'sd2213}, {9'sd-182, 13'sd2233, 13'sd-2107}},
{{11'sd837, 13'sd2533, 13'sd3136}, {10'sd422, 10'sd345, 12'sd1908}, {11'sd-990, 11'sd-786, 13'sd2569}},
{{12'sd-1104, 12'sd-1364, 11'sd663}, {10'sd-367, 13'sd-2208, 13'sd2399}, {13'sd2575, 12'sd1057, 12'sd-1138}},
{{11'sd-703, 11'sd-871, 12'sd1644}, {10'sd409, 13'sd-3472, 12'sd-1640}, {10'sd480, 12'sd-1848, 11'sd726}},
{{13'sd-2923, 12'sd-1229, 13'sd3013}, {12'sd-1699, 13'sd-2330, 11'sd-647}, {12'sd-1208, 13'sd2135, 9'sd-161}},
{{13'sd2512, 11'sd793, 12'sd-1508}, {13'sd3557, 13'sd2448, 12'sd1299}, {13'sd2199, 13'sd2854, 12'sd-1288}},
{{11'sd842, 10'sd453, 13'sd-2977}, {11'sd724, 11'sd-684, 13'sd-2260}, {6'sd-30, 12'sd-1652, 12'sd-1791}},
{{11'sd972, 13'sd2382, 13'sd2573}, {12'sd-1879, 11'sd-684, 9'sd-205}, {13'sd2779, 11'sd573, 11'sd669}},
{{11'sd894, 12'sd1827, 11'sd953}, {12'sd-1809, 9'sd-210, 13'sd-3037}, {12'sd1518, 11'sd-754, 12'sd1249}},
{{13'sd2250, 12'sd-1713, 12'sd1397}, {12'sd-1402, 12'sd2012, 12'sd-1283}, {11'sd-919, 13'sd2278, 13'sd2221}},
{{4'sd7, 12'sd-1242, 10'sd-332}, {14'sd-4212, 10'sd285, 12'sd1284}, {12'sd-1166, 13'sd-3112, 12'sd-1960}},
{{12'sd-1439, 12'sd1764, 12'sd2031}, {13'sd2483, 8'sd79, 13'sd2342}, {12'sd2046, 13'sd2457, 12'sd1965}},
{{13'sd-3128, 13'sd-2178, 13'sd-3793}, {12'sd-1255, 11'sd-815, 11'sd788}, {11'sd-864, 13'sd-2407, 13'sd-2512}},
{{13'sd-2857, 13'sd-2992, 8'sd94}, {12'sd1028, 9'sd-229, 12'sd-1249}, {12'sd1152, 12'sd1719, 12'sd-1758}},
{{12'sd-1337, 13'sd-2404, 7'sd-54}, {13'sd-3103, 12'sd-1402, 9'sd-252}, {10'sd-347, 13'sd-2573, 12'sd1410}},
{{13'sd-2453, 12'sd1475, 11'sd955}, {12'sd-1978, 8'sd119, 11'sd753}, {13'sd-2625, 12'sd1368, 13'sd-2666}},
{{12'sd1525, 13'sd2359, 13'sd-2570}, {11'sd-913, 12'sd-1373, 12'sd-1835}, {13'sd2222, 12'sd-1519, 11'sd619}},
{{10'sd-261, 11'sd554, 11'sd-923}, {9'sd-225, 12'sd-1031, 13'sd-2485}, {13'sd-2433, 13'sd-2385, 11'sd578}},
{{13'sd2370, 13'sd3183, 12'sd-1715}, {12'sd-1137, 11'sd-802, 12'sd-1673}, {13'sd2347, 13'sd-2117, 13'sd2713}},
{{11'sd-1004, 12'sd-1563, 11'sd900}, {13'sd3301, 12'sd1491, 11'sd981}, {11'sd-790, 11'sd-817, 12'sd-1476}}},
{
{{10'sd-390, 12'sd1186, 12'sd1695}, {12'sd-1571, 11'sd-549, 12'sd-1335}, {7'sd-62, 11'sd655, 12'sd-1442}},
{{11'sd-581, 12'sd1358, 9'sd-221}, {12'sd1068, 10'sd455, 8'sd121}, {9'sd141, 6'sd31, 12'sd-1978}},
{{12'sd1750, 13'sd2363, 12'sd-1900}, {11'sd964, 11'sd-618, 11'sd-728}, {12'sd-1098, 12'sd1554, 12'sd-1182}},
{{12'sd1114, 10'sd-475, 12'sd1063}, {11'sd590, 11'sd529, 10'sd-329}, {12'sd-1584, 13'sd-2220, 9'sd152}},
{{11'sd683, 13'sd-3430, 13'sd-2942}, {13'sd-2569, 9'sd239, 8'sd-87}, {13'sd-2437, 10'sd481, 12'sd-1127}},
{{13'sd-2371, 12'sd1116, 13'sd3855}, {11'sd571, 12'sd-1379, 13'sd2261}, {12'sd-1771, 12'sd-1359, 12'sd1999}},
{{7'sd-45, 8'sd-83, 11'sd679}, {12'sd-1714, 11'sd895, 5'sd-10}, {12'sd1783, 12'sd-1832, 13'sd2957}},
{{13'sd2149, 13'sd2884, 13'sd-2309}, {11'sd-695, 13'sd2061, 13'sd2574}, {13'sd2543, 12'sd1624, 12'sd-1980}},
{{12'sd-1856, 10'sd-359, 12'sd-1229}, {13'sd-2876, 13'sd-2976, 13'sd-2914}, {12'sd1189, 11'sd-829, 10'sd322}},
{{9'sd-175, 13'sd-2091, 8'sd72}, {12'sd-1324, 12'sd-1580, 8'sd103}, {9'sd253, 13'sd2087, 13'sd-2381}},
{{8'sd-104, 13'sd-2270, 6'sd22}, {13'sd-2526, 9'sd236, 12'sd-1356}, {12'sd-1547, 11'sd-630, 13'sd2392}},
{{11'sd620, 11'sd-522, 12'sd-1878}, {11'sd-836, 12'sd1175, 13'sd-2086}, {12'sd-1775, 13'sd2198, 10'sd451}},
{{13'sd-2278, 12'sd-1102, 13'sd-2759}, {11'sd-713, 6'sd-28, 12'sd-1548}, {13'sd-2860, 12'sd-2029, 12'sd1574}},
{{11'sd-994, 12'sd2005, 13'sd-2149}, {13'sd-2587, 10'sd-301, 13'sd-2550}, {12'sd-1876, 10'sd453, 13'sd-2558}},
{{11'sd-647, 8'sd89, 11'sd799}, {13'sd-3741, 13'sd-2502, 13'sd2290}, {12'sd1456, 12'sd-1990, 12'sd-1032}},
{{11'sd-762, 13'sd-2511, 11'sd792}, {11'sd-883, 13'sd-3201, 11'sd-997}, {10'sd444, 12'sd1518, 12'sd-1890}},
{{11'sd-665, 12'sd-1236, 9'sd201}, {13'sd2144, 10'sd306, 13'sd2389}, {11'sd-616, 10'sd-444, 12'sd-1579}},
{{12'sd-1376, 11'sd-1007, 12'sd1707}, {13'sd-2989, 12'sd1454, 13'sd-2375}, {13'sd-3363, 12'sd1788, 11'sd-715}},
{{12'sd-1255, 11'sd-950, 12'sd-1891}, {12'sd-1109, 10'sd291, 12'sd1977}, {13'sd2635, 13'sd2212, 12'sd1131}},
{{12'sd1194, 12'sd1700, 13'sd2883}, {10'sd388, 9'sd205, 12'sd1973}, {13'sd2223, 5'sd13, 12'sd-1156}},
{{13'sd2618, 12'sd-1230, 1'sd0}, {8'sd75, 6'sd-19, 10'sd435}, {10'sd337, 12'sd1671, 11'sd962}},
{{12'sd1347, 12'sd1951, 12'sd-1793}, {9'sd-176, 11'sd-880, 13'sd2096}, {12'sd-1753, 12'sd1459, 11'sd-873}},
{{12'sd-1791, 10'sd509, 10'sd455}, {9'sd194, 13'sd-2541, 13'sd-2401}, {13'sd2125, 13'sd-2737, 11'sd537}},
{{11'sd-623, 12'sd1659, 10'sd-256}, {12'sd-1072, 12'sd-1694, 11'sd-964}, {12'sd1941, 12'sd1090, 13'sd2398}},
{{13'sd-2526, 12'sd1921, 13'sd2070}, {12'sd1089, 11'sd963, 12'sd-1545}, {12'sd1129, 13'sd-2592, 13'sd-2453}},
{{12'sd1306, 12'sd1069, 11'sd-605}, {11'sd-1021, 11'sd-986, 12'sd-1239}, {12'sd-1759, 11'sd-586, 11'sd739}},
{{12'sd-1252, 12'sd-1188, 13'sd2234}, {10'sd-400, 12'sd-1494, 9'sd-179}, {12'sd1163, 11'sd-827, 13'sd2336}},
{{10'sd458, 13'sd-2827, 12'sd1969}, {11'sd-790, 9'sd128, 8'sd64}, {13'sd-2219, 12'sd2003, 13'sd2129}},
{{12'sd-1066, 13'sd2923, 9'sd-132}, {10'sd-372, 13'sd2087, 12'sd1619}, {12'sd-1669, 12'sd1575, 13'sd2106}},
{{13'sd-2127, 9'sd173, 8'sd83}, {12'sd-1107, 6'sd20, 12'sd-2010}, {11'sd-545, 9'sd-229, 12'sd-1402}},
{{13'sd-2213, 13'sd-2444, 13'sd-2079}, {13'sd2395, 11'sd514, 11'sd-645}, {12'sd-1464, 5'sd11, 13'sd-2417}},
{{13'sd2519, 13'sd-2285, 12'sd-1300}, {10'sd-442, 13'sd-2613, 13'sd2202}, {8'sd-123, 8'sd-79, 13'sd2851}},
{{7'sd50, 12'sd-1477, 12'sd-1316}, {12'sd1942, 13'sd2741, 10'sd489}, {11'sd-703, 13'sd2566, 12'sd1406}},
{{11'sd-1017, 12'sd-1548, 12'sd1513}, {11'sd-817, 7'sd37, 12'sd-1947}, {7'sd40, 12'sd-1474, 12'sd-1775}},
{{10'sd268, 12'sd1434, 12'sd1940}, {13'sd2939, 10'sd-438, 12'sd-1958}, {11'sd564, 12'sd1264, 10'sd-414}},
{{13'sd2170, 11'sd-956, 9'sd-189}, {11'sd-880, 13'sd-2484, 12'sd1924}, {8'sd-108, 13'sd-2262, 12'sd-1405}},
{{11'sd596, 12'sd1703, 10'sd-283}, {10'sd-258, 9'sd-221, 12'sd1810}, {11'sd-1014, 10'sd311, 13'sd3061}},
{{11'sd709, 12'sd1708, 12'sd1104}, {11'sd-566, 13'sd-2636, 11'sd-963}, {10'sd275, 13'sd-2121, 12'sd1533}},
{{6'sd29, 12'sd1964, 13'sd2835}, {12'sd1233, 12'sd1694, 11'sd-923}, {10'sd502, 4'sd-4, 7'sd-46}},
{{12'sd1740, 13'sd2461, 12'sd-1224}, {10'sd271, 12'sd1200, 11'sd-926}, {11'sd767, 13'sd2128, 11'sd-531}},
{{10'sd262, 12'sd1307, 12'sd-2035}, {13'sd-2342, 9'sd182, 11'sd-802}, {13'sd-3265, 10'sd-388, 12'sd1030}},
{{13'sd-2271, 12'sd-1291, 12'sd1853}, {13'sd-2899, 13'sd-3139, 12'sd-1532}, {12'sd-1374, 12'sd1671, 12'sd1671}},
{{10'sd388, 13'sd2713, 13'sd2768}, {8'sd-122, 13'sd2794, 13'sd-2088}, {13'sd-2370, 12'sd-1176, 13'sd2139}},
{{13'sd2663, 13'sd2796, 13'sd3424}, {10'sd463, 11'sd-702, 12'sd2031}, {13'sd-3105, 12'sd-1287, 13'sd-2638}},
{{13'sd-2753, 13'sd2400, 12'sd-1045}, {13'sd2296, 7'sd46, 11'sd792}, {10'sd402, 12'sd-1719, 12'sd-1232}},
{{12'sd2006, 13'sd2718, 11'sd-637}, {12'sd-1154, 12'sd1795, 9'sd181}, {12'sd-1169, 12'sd1455, 11'sd776}},
{{11'sd-818, 12'sd1533, 9'sd177}, {11'sd864, 11'sd529, 11'sd773}, {10'sd380, 12'sd1362, 7'sd33}},
{{12'sd-1619, 12'sd1382, 12'sd1615}, {12'sd1626, 8'sd-102, 10'sd-423}, {11'sd680, 10'sd-462, 12'sd2025}},
{{11'sd-592, 13'sd2766, 9'sd242}, {13'sd-2317, 12'sd1075, 12'sd1858}, {12'sd-1499, 11'sd-976, 13'sd3170}},
{{11'sd828, 13'sd-2337, 13'sd2152}, {11'sd761, 12'sd-1380, 12'sd-1280}, {13'sd-2153, 13'sd2737, 12'sd-1291}},
{{12'sd-1684, 9'sd218, 13'sd2116}, {9'sd236, 13'sd-2289, 12'sd1831}, {12'sd1432, 11'sd-940, 11'sd-916}},
{{11'sd662, 13'sd2066, 13'sd-2054}, {11'sd-679, 10'sd-448, 12'sd1769}, {11'sd-688, 11'sd-695, 12'sd1121}},
{{11'sd-778, 9'sd-179, 10'sd466}, {13'sd2605, 12'sd1662, 10'sd-452}, {13'sd-2215, 12'sd2007, 12'sd-1883}},
{{13'sd2298, 11'sd-554, 11'sd-997}, {12'sd-1328, 11'sd-820, 12'sd-2038}, {11'sd-723, 4'sd4, 12'sd-1251}},
{{13'sd-2323, 12'sd-1331, 12'sd-1547}, {11'sd-787, 11'sd-623, 11'sd-800}, {13'sd-2796, 12'sd-2016, 12'sd1114}},
{{12'sd-1462, 12'sd-1449, 13'sd-2239}, {12'sd1094, 10'sd352, 12'sd2035}, {13'sd2896, 13'sd3320, 12'sd-1732}},
{{11'sd685, 13'sd-3582, 10'sd-311}, {14'sd-4259, 12'sd-1686, 12'sd-1068}, {13'sd-2907, 13'sd-3526, 12'sd-1398}},
{{9'sd-141, 10'sd299, 9'sd-217}, {11'sd-753, 10'sd-452, 11'sd-946}, {13'sd-3221, 11'sd-728, 9'sd-132}},
{{11'sd-966, 11'sd868, 11'sd-978}, {11'sd-513, 12'sd-1811, 12'sd1774}, {12'sd1508, 12'sd1562, 11'sd872}},
{{12'sd1244, 10'sd-261, 12'sd1273}, {11'sd557, 12'sd-1117, 12'sd1509}, {11'sd955, 12'sd-1615, 12'sd1431}},
{{12'sd-1510, 13'sd2676, 12'sd2040}, {10'sd390, 10'sd-438, 13'sd-2409}, {13'sd-2553, 12'sd1995, 12'sd-1158}},
{{13'sd-2150, 13'sd2233, 13'sd-2705}, {10'sd-486, 11'sd882, 13'sd-2903}, {12'sd1746, 12'sd1554, 12'sd-1070}},
{{9'sd-146, 12'sd1482, 11'sd-939}, {13'sd2455, 12'sd1073, 13'sd2329}, {13'sd-2644, 12'sd-2032, 9'sd-143}},
{{12'sd1463, 13'sd2622, 13'sd2123}, {13'sd2551, 12'sd1520, 12'sd1187}, {11'sd-777, 12'sd1364, 12'sd2045}}},
{
{{13'sd-2331, 11'sd-577, 13'sd-2334}, {10'sd282, 13'sd-2396, 12'sd-1196}, {13'sd2292, 12'sd2046, 12'sd1996}},
{{10'sd-325, 13'sd-2224, 13'sd-2777}, {12'sd1469, 11'sd-903, 11'sd-715}, {12'sd-1756, 13'sd-2214, 10'sd423}},
{{9'sd208, 12'sd-1638, 12'sd1499}, {11'sd540, 10'sd-445, 9'sd-187}, {10'sd267, 13'sd2519, 13'sd2760}},
{{12'sd1866, 13'sd2307, 13'sd-2052}, {12'sd1311, 10'sd-449, 13'sd2184}, {12'sd-1318, 12'sd1525, 12'sd-1923}},
{{13'sd-2474, 14'sd-4254, 13'sd-3460}, {10'sd445, 9'sd-132, 13'sd-3987}, {13'sd3769, 13'sd3747, 12'sd-1575}},
{{12'sd-1478, 14'sd-4749, 12'sd1672}, {13'sd-3410, 13'sd-3184, 13'sd-2959}, {11'sd-739, 12'sd1707, 10'sd-334}},
{{11'sd633, 12'sd-1555, 13'sd2771}, {13'sd-2724, 13'sd-3728, 12'sd-1800}, {12'sd-1029, 12'sd-1706, 12'sd2036}},
{{12'sd1699, 12'sd1478, 11'sd-986}, {13'sd2155, 12'sd-1964, 13'sd2109}, {11'sd-579, 11'sd928, 12'sd-1579}},
{{13'sd-2838, 12'sd-1309, 12'sd-2047}, {12'sd-1870, 10'sd-432, 13'sd-2713}, {9'sd-204, 9'sd251, 12'sd-1387}},
{{13'sd3609, 13'sd2943, 12'sd1749}, {11'sd-1008, 13'sd2139, 11'sd833}, {12'sd1159, 13'sd3182, 9'sd-234}},
{{12'sd1735, 11'sd-577, 13'sd-2423}, {11'sd-723, 12'sd1027, 13'sd-3215}, {13'sd2970, 12'sd1655, 12'sd1091}},
{{12'sd-1054, 9'sd242, 5'sd11}, {11'sd513, 13'sd2220, 13'sd-2524}, {13'sd-2121, 12'sd-1118, 12'sd-1347}},
{{13'sd3214, 12'sd1615, 13'sd-3430}, {10'sd-467, 13'sd-2371, 13'sd-2664}, {13'sd3187, 14'sd4237, 13'sd2948}},
{{13'sd2608, 10'sd328, 12'sd-1372}, {12'sd1573, 9'sd225, 12'sd-1100}, {12'sd-1538, 12'sd1445, 11'sd-527}},
{{14'sd-4395, 7'sd45, 11'sd-851}, {13'sd3011, 12'sd1818, 13'sd2409}, {12'sd1405, 8'sd65, 12'sd1734}},
{{11'sd773, 12'sd1730, 11'sd-895}, {12'sd-1211, 13'sd-2253, 13'sd-2696}, {9'sd-218, 10'sd351, 11'sd794}},
{{11'sd795, 7'sd38, 13'sd2457}, {10'sd378, 13'sd-2305, 12'sd-1275}, {8'sd107, 12'sd-1324, 12'sd-1511}},
{{13'sd-2857, 13'sd-2588, 12'sd-1916}, {11'sd-760, 11'sd-740, 12'sd-1934}, {13'sd2050, 8'sd-65, 10'sd-336}},
{{13'sd2355, 11'sd-787, 12'sd-1528}, {9'sd232, 13'sd2256, 12'sd-2023}, {12'sd1626, 12'sd1877, 11'sd794}},
{{13'sd2213, 12'sd-1729, 13'sd3559}, {13'sd-2599, 12'sd1595, 13'sd2795}, {12'sd-1996, 12'sd-2023, 11'sd916}},
{{13'sd-2569, 12'sd-1570, 11'sd-823}, {12'sd-1697, 12'sd1739, 12'sd-1665}, {11'sd-533, 11'sd-546, 12'sd1658}},
{{12'sd-1868, 11'sd-673, 9'sd142}, {11'sd-554, 10'sd461, 13'sd2803}, {13'sd-2638, 11'sd925, 12'sd-2032}},
{{13'sd2830, 11'sd-1011, 12'sd1979}, {10'sd-435, 9'sd201, 12'sd1349}, {11'sd-773, 11'sd809, 11'sd698}},
{{13'sd2055, 10'sd446, 12'sd-1288}, {13'sd-2688, 13'sd3147, 10'sd447}, {11'sd-801, 13'sd-2621, 12'sd-1480}},
{{9'sd188, 13'sd3009, 12'sd-1177}, {12'sd-1736, 12'sd1136, 12'sd-1838}, {12'sd1440, 9'sd216, 12'sd-1805}},
{{11'sd760, 12'sd-1327, 13'sd-3510}, {13'sd3176, 12'sd1418, 12'sd1484}, {12'sd1611, 13'sd2508, 12'sd1508}},
{{9'sd219, 13'sd-2160, 14'sd-4409}, {12'sd-2010, 13'sd-2701, 14'sd-4941}, {14'sd-4854, 10'sd-340, 12'sd-1567}},
{{12'sd-2035, 9'sd-136, 13'sd-2338}, {13'sd-2711, 9'sd-219, 10'sd466}, {12'sd-1187, 12'sd1339, 12'sd1949}},
{{11'sd587, 12'sd1090, 12'sd1343}, {12'sd1035, 12'sd-1455, 13'sd2990}, {13'sd2341, 12'sd1263, 10'sd-340}},
{{13'sd-2399, 13'sd2320, 9'sd234}, {13'sd-3547, 9'sd-223, 13'sd-3278}, {10'sd464, 4'sd4, 9'sd-248}},
{{13'sd2693, 13'sd2918, 13'sd-2344}, {13'sd2552, 11'sd793, 12'sd-1624}, {12'sd-1971, 12'sd-1036, 12'sd1581}},
{{13'sd-2394, 12'sd-1905, 13'sd2240}, {12'sd2047, 12'sd-1318, 11'sd-719}, {13'sd2224, 13'sd2617, 12'sd1529}},
{{13'sd-2108, 12'sd-2020, 12'sd1167}, {12'sd-1549, 13'sd-2286, 10'sd391}, {13'sd-3668, 12'sd1301, 12'sd-1891}},
{{12'sd1965, 12'sd-1712, 10'sd-456}, {12'sd1558, 12'sd1730, 12'sd-1933}, {11'sd795, 11'sd532, 13'sd-2473}},
{{13'sd-2656, 10'sd-320, 10'sd-510}, {13'sd-2129, 13'sd2746, 12'sd1709}, {12'sd-1504, 12'sd1651, 6'sd23}},
{{11'sd-557, 11'sd882, 11'sd558}, {12'sd1567, 12'sd-1941, 13'sd2283}, {11'sd580, 13'sd-2460, 12'sd-1408}},
{{11'sd-916, 12'sd-1205, 13'sd3116}, {11'sd-548, 13'sd-3540, 10'sd266}, {14'sd-4935, 12'sd-1394, 11'sd-767}},
{{10'sd-269, 13'sd-2805, 13'sd-3938}, {12'sd-1118, 12'sd-1284, 11'sd-806}, {11'sd-638, 11'sd-879, 13'sd-2353}},
{{11'sd-597, 13'sd-2250, 11'sd945}, {13'sd-2082, 10'sd-269, 12'sd1542}, {12'sd-1273, 13'sd2398, 12'sd1534}},
{{13'sd-2803, 11'sd-996, 12'sd1531}, {11'sd-711, 13'sd2160, 12'sd-1778}, {12'sd-1240, 11'sd-831, 12'sd-1829}},
{{11'sd-819, 11'sd753, 12'sd1061}, {13'sd-2255, 13'sd-2366, 12'sd-1354}, {14'sd-4150, 13'sd-2609, 13'sd-3446}},
{{9'sd-141, 13'sd-2248, 12'sd-1041}, {12'sd1452, 10'sd385, 12'sd-1083}, {13'sd3227, 14'sd5794, 14'sd4938}},
{{11'sd1011, 9'sd-142, 12'sd-1803}, {13'sd-2304, 13'sd2499, 11'sd-797}, {12'sd1523, 14'sd5442, 13'sd3937}},
{{13'sd3776, 13'sd-2697, 14'sd-5309}, {8'sd-73, 14'sd-7208, 13'sd-2785}, {12'sd1675, 10'sd-447, 13'sd-2959}},
{{12'sd-1186, 13'sd-2598, 13'sd-2239}, {12'sd-1524, 11'sd550, 10'sd-298}, {12'sd1463, 12'sd1410, 13'sd-2088}},
{{13'sd-2454, 12'sd1686, 11'sd873}, {13'sd-3335, 11'sd-704, 6'sd19}, {11'sd-786, 9'sd252, 9'sd-198}},
{{13'sd-3396, 12'sd1700, 12'sd1147}, {12'sd-1511, 11'sd864, 12'sd-1376}, {14'sd-4861, 13'sd-2397, 12'sd1054}},
{{9'sd234, 12'sd-1533, 13'sd-2394}, {13'sd-3524, 11'sd522, 13'sd-3280}, {11'sd666, 12'sd1641, 13'sd-2936}},
{{10'sd259, 11'sd537, 13'sd-2339}, {12'sd1336, 11'sd542, 12'sd1356}, {12'sd-1078, 13'sd-2658, 12'sd1531}},
{{11'sd-665, 12'sd1999, 13'sd3249}, {12'sd1957, 11'sd826, 12'sd1980}, {13'sd-2685, 12'sd1904, 12'sd-1799}},
{{10'sd-409, 11'sd665, 10'sd-478}, {12'sd1284, 11'sd-1019, 11'sd654}, {12'sd1695, 13'sd2620, 12'sd1472}},
{{13'sd3470, 12'sd-1167, 13'sd-2330}, {12'sd1833, 10'sd453, 12'sd-1524}, {14'sd4682, 10'sd-327, 13'sd2297}},
{{8'sd-76, 10'sd-382, 6'sd-16}, {12'sd1661, 9'sd-149, 11'sd898}, {14'sd6343, 14'sd4315, 13'sd2829}},
{{11'sd-961, 13'sd-2736, 13'sd2675}, {13'sd-3009, 13'sd-2982, 9'sd-178}, {13'sd-2453, 12'sd1937, 12'sd-1245}},
{{9'sd179, 9'sd-174, 14'sd-5158}, {13'sd2537, 12'sd-1862, 12'sd-1948}, {13'sd-2055, 10'sd313, 13'sd2919}},
{{12'sd-1690, 11'sd913, 13'sd3724}, {12'sd-1726, 13'sd2149, 12'sd1197}, {13'sd-2606, 13'sd-2429, 7'sd58}},
{{11'sd-745, 13'sd2296, 14'sd-4614}, {12'sd-1930, 12'sd-1169, 10'sd323}, {14'sd8089, 14'sd4791, 12'sd1080}},
{{11'sd-576, 13'sd-2362, 12'sd-1317}, {11'sd-566, 11'sd-736, 12'sd1211}, {9'sd-236, 12'sd-1243, 11'sd718}},
{{12'sd-1771, 12'sd1579, 12'sd1111}, {12'sd1288, 12'sd-1587, 13'sd-2500}, {13'sd2867, 12'sd-1285, 12'sd1885}},
{{8'sd-102, 12'sd-2000, 12'sd-1438}, {11'sd719, 12'sd-1430, 12'sd-1370}, {14'sd-5216, 13'sd-3028, 13'sd-3383}},
{{13'sd-3376, 12'sd-1101, 8'sd116}, {11'sd-994, 13'sd2060, 11'sd780}, {12'sd-1616, 10'sd336, 12'sd1323}},
{{11'sd957, 13'sd-2626, 12'sd-1184}, {11'sd-920, 10'sd273, 11'sd-549}, {13'sd3619, 12'sd-1251, 12'sd1902}},
{{11'sd828, 10'sd444, 10'sd286}, {13'sd-2066, 13'sd-3173, 12'sd1914}, {12'sd-1282, 11'sd-762, 12'sd-1645}},
{{11'sd892, 8'sd91, 13'sd2381}, {13'sd3944, 7'sd61, 13'sd3646}, {11'sd778, 11'sd-904, 12'sd1786}}},
{
{{12'sd1151, 12'sd1356, 11'sd-557}, {11'sd1012, 12'sd-1536, 12'sd-1319}, {11'sd776, 13'sd2223, 10'sd268}},
{{13'sd-2890, 11'sd933, 13'sd-2181}, {13'sd-2650, 12'sd1255, 11'sd1008}, {11'sd-882, 12'sd-1512, 13'sd2442}},
{{12'sd-1678, 12'sd1619, 12'sd1264}, {11'sd980, 7'sd-48, 11'sd-629}, {12'sd1768, 10'sd358, 13'sd2244}},
{{8'sd-101, 9'sd133, 12'sd1132}, {13'sd-2323, 12'sd-1039, 12'sd-1334}, {13'sd-2075, 10'sd336, 7'sd-39}},
{{10'sd-417, 12'sd1311, 12'sd1352}, {12'sd-1564, 11'sd669, 12'sd1678}, {12'sd-1513, 13'sd2908, 13'sd2594}},
{{10'sd316, 12'sd-1704, 10'sd-343}, {10'sd-479, 10'sd468, 12'sd-1438}, {10'sd-266, 9'sd208, 13'sd2298}},
{{10'sd287, 10'sd-401, 8'sd126}, {13'sd2141, 12'sd-1802, 12'sd1973}, {12'sd1778, 12'sd1279, 12'sd-1551}},
{{12'sd-1758, 9'sd211, 11'sd654}, {12'sd1747, 2'sd-1, 13'sd-2402}, {12'sd-1313, 11'sd697, 11'sd622}},
{{12'sd-1587, 11'sd-899, 12'sd1458}, {11'sd937, 12'sd-2010, 11'sd951}, {12'sd2001, 13'sd2687, 12'sd-1181}},
{{9'sd-228, 12'sd-1983, 12'sd1302}, {10'sd-270, 13'sd2735, 10'sd273}, {11'sd860, 12'sd1334, 12'sd-2046}},
{{12'sd1391, 10'sd-497, 12'sd1980}, {13'sd2235, 12'sd-1672, 10'sd-454}, {12'sd1646, 10'sd488, 10'sd-471}},
{{13'sd2066, 13'sd2230, 9'sd135}, {10'sd449, 12'sd1462, 13'sd-2417}, {11'sd733, 12'sd1809, 13'sd2399}},
{{13'sd-2552, 12'sd1120, 13'sd2283}, {13'sd-2406, 12'sd-1259, 13'sd2763}, {12'sd-1458, 12'sd1273, 8'sd-124}},
{{13'sd-2496, 8'sd-96, 12'sd-1340}, {11'sd914, 11'sd-722, 13'sd-2756}, {10'sd-459, 13'sd-2662, 9'sd227}},
{{13'sd2733, 11'sd838, 12'sd-1345}, {12'sd-1267, 9'sd233, 13'sd2168}, {11'sd-940, 12'sd1239, 13'sd2497}},
{{12'sd1361, 13'sd2181, 13'sd2809}, {12'sd-1358, 13'sd2431, 13'sd2157}, {13'sd-2775, 11'sd836, 7'sd46}},
{{11'sd1000, 10'sd396, 12'sd-1610}, {12'sd-2037, 12'sd-1896, 10'sd-458}, {12'sd1117, 11'sd889, 11'sd-580}},
{{11'sd842, 12'sd1359, 13'sd2617}, {13'sd2138, 13'sd-2640, 13'sd-2058}, {12'sd1981, 13'sd2422, 12'sd1982}},
{{13'sd-2158, 9'sd154, 12'sd1119}, {11'sd573, 12'sd-1578, 12'sd-2041}, {13'sd2557, 10'sd-440, 10'sd428}},
{{12'sd1619, 10'sd-301, 11'sd652}, {13'sd2598, 13'sd2479, 11'sd-691}, {13'sd2811, 13'sd2684, 13'sd2295}},
{{9'sd148, 9'sd-150, 12'sd1466}, {13'sd-2531, 11'sd-995, 13'sd2475}, {12'sd-1709, 11'sd949, 13'sd2324}},
{{9'sd-196, 12'sd1673, 13'sd2728}, {11'sd-588, 11'sd658, 12'sd-1328}, {12'sd1793, 12'sd1562, 11'sd-541}},
{{12'sd1628, 6'sd-16, 11'sd-515}, {11'sd-851, 12'sd-1853, 13'sd-2358}, {10'sd467, 12'sd-1702, 12'sd-1332}},
{{4'sd5, 12'sd-1928, 13'sd2703}, {13'sd2545, 10'sd-447, 11'sd878}, {12'sd1259, 12'sd-1769, 12'sd1177}},
{{9'sd-190, 10'sd-445, 10'sd-275}, {13'sd2597, 10'sd314, 12'sd1106}, {13'sd-2165, 12'sd-1443, 13'sd2111}},
{{13'sd2249, 9'sd-143, 8'sd-115}, {12'sd1038, 12'sd-1261, 12'sd2045}, {12'sd-1699, 11'sd-1018, 9'sd-184}},
{{13'sd-2586, 13'sd2698, 12'sd1634}, {13'sd-2060, 10'sd-327, 13'sd-3571}, {10'sd-422, 13'sd-2775, 10'sd-483}},
{{13'sd2191, 13'sd2564, 9'sd165}, {11'sd680, 13'sd2726, 12'sd1740}, {12'sd1266, 12'sd-1199, 12'sd1727}},
{{13'sd2051, 12'sd1235, 12'sd1699}, {12'sd-1344, 8'sd68, 13'sd-2524}, {11'sd-801, 11'sd-590, 13'sd-2453}},
{{13'sd-2259, 12'sd1589, 9'sd224}, {10'sd-494, 10'sd306, 13'sd2629}, {13'sd2536, 11'sd-738, 12'sd1213}},
{{10'sd375, 13'sd2600, 10'sd306}, {13'sd-2321, 11'sd-562, 12'sd-1717}, {10'sd343, 11'sd-734, 13'sd2079}},
{{12'sd-1783, 12'sd-1377, 9'sd184}, {11'sd765, 11'sd773, 12'sd1805}, {11'sd863, 12'sd1657, 10'sd320}},
{{8'sd-68, 11'sd-696, 9'sd-180}, {11'sd-656, 11'sd-869, 12'sd1373}, {12'sd-1140, 12'sd1835, 10'sd-394}},
{{10'sd-309, 10'sd-466, 12'sd-1421}, {11'sd-637, 12'sd-2020, 10'sd416}, {11'sd-893, 13'sd-2381, 12'sd1530}},
{{13'sd2074, 12'sd1517, 12'sd1346}, {13'sd2617, 9'sd154, 13'sd-2691}, {8'sd117, 13'sd2084, 11'sd701}},
{{9'sd-237, 13'sd2421, 12'sd2047}, {11'sd-1019, 13'sd-2722, 13'sd2180}, {12'sd-1845, 10'sd354, 13'sd-2325}},
{{12'sd-1713, 11'sd602, 9'sd201}, {11'sd546, 11'sd921, 13'sd-3027}, {12'sd1643, 13'sd2940, 12'sd-1811}},
{{12'sd-1031, 11'sd-610, 12'sd-1347}, {12'sd-1500, 12'sd1932, 12'sd1312}, {12'sd1191, 12'sd1571, 11'sd-973}},
{{13'sd2520, 13'sd2171, 6'sd-22}, {12'sd1975, 12'sd-1060, 13'sd2467}, {11'sd-818, 12'sd-1297, 12'sd1791}},
{{8'sd105, 11'sd-680, 13'sd-2116}, {12'sd-1476, 13'sd-2614, 13'sd-2524}, {12'sd-1539, 8'sd66, 10'sd-495}},
{{10'sd383, 12'sd-1510, 12'sd1786}, {12'sd1763, 13'sd2365, 13'sd2685}, {11'sd976, 12'sd1531, 10'sd-389}},
{{12'sd1538, 11'sd828, 11'sd-625}, {12'sd-1434, 12'sd-1321, 12'sd1353}, {13'sd2082, 7'sd60, 11'sd723}},
{{12'sd-1342, 11'sd928, 12'sd1181}, {11'sd-1022, 10'sd-505, 11'sd-515}, {12'sd-1963, 13'sd-2334, 11'sd885}},
{{14'sd-4136, 13'sd-2649, 8'sd-127}, {13'sd-3387, 11'sd-660, 9'sd-189}, {12'sd-1518, 11'sd931, 12'sd-1861}},
{{11'sd-795, 12'sd1643, 12'sd1728}, {13'sd2499, 10'sd285, 13'sd-2606}, {11'sd-711, 12'sd1402, 12'sd-1626}},
{{12'sd1425, 8'sd72, 10'sd-309}, {12'sd-1203, 11'sd1001, 7'sd-56}, {9'sd165, 12'sd-1403, 12'sd1384}},
{{13'sd2602, 10'sd509, 13'sd-2194}, {9'sd-248, 11'sd-608, 13'sd2164}, {12'sd1097, 13'sd-2279, 11'sd-725}},
{{10'sd-301, 13'sd2422, 12'sd-1443}, {11'sd-901, 13'sd2457, 13'sd-2688}, {12'sd1187, 13'sd2417, 12'sd1677}},
{{12'sd-1165, 13'sd-2381, 12'sd-1502}, {11'sd966, 13'sd-2137, 12'sd2016}, {10'sd453, 11'sd807, 11'sd-825}},
{{12'sd1800, 11'sd-619, 13'sd2102}, {9'sd203, 12'sd1832, 13'sd-2552}, {12'sd-1949, 13'sd2596, 13'sd-3217}},
{{13'sd2257, 13'sd2620, 13'sd2090}, {11'sd967, 11'sd776, 12'sd1749}, {13'sd2329, 12'sd1431, 9'sd211}},
{{11'sd737, 12'sd-1093, 12'sd-1954}, {9'sd-199, 13'sd2433, 11'sd-760}, {7'sd52, 5'sd9, 12'sd1442}},
{{10'sd-433, 9'sd-180, 12'sd-1538}, {10'sd257, 5'sd-13, 13'sd2411}, {12'sd-1599, 13'sd-3079, 12'sd1533}},
{{13'sd2132, 13'sd-2427, 13'sd2586}, {12'sd-1171, 13'sd-2573, 12'sd-1274}, {13'sd2408, 12'sd1262, 11'sd811}},
{{11'sd-836, 10'sd-360, 10'sd-409}, {12'sd-1664, 11'sd783, 12'sd1488}, {12'sd1549, 12'sd1061, 13'sd2329}},
{{11'sd-677, 13'sd-2433, 12'sd-1506}, {13'sd2346, 10'sd357, 11'sd-540}, {13'sd-2290, 4'sd-7, 12'sd1803}},
{{10'sd445, 12'sd-1132, 13'sd2522}, {13'sd2590, 12'sd1906, 13'sd2396}, {12'sd1055, 12'sd1853, 13'sd3579}},
{{12'sd1111, 13'sd3138, 10'sd447}, {12'sd1051, 10'sd413, 9'sd227}, {11'sd580, 13'sd-2802, 12'sd-1164}},
{{13'sd2694, 8'sd-101, 12'sd1031}, {12'sd-1189, 12'sd1799, 8'sd-123}, {12'sd-1482, 13'sd2519, 11'sd-974}},
{{13'sd2881, 13'sd2085, 12'sd-1394}, {11'sd519, 11'sd-848, 12'sd1308}, {13'sd2966, 12'sd1980, 12'sd1092}},
{{11'sd959, 12'sd1581, 13'sd2728}, {12'sd-1822, 13'sd-2500, 10'sd-303}, {12'sd-1291, 12'sd1956, 12'sd-1183}},
{{13'sd-2204, 13'sd2388, 10'sd283}, {12'sd1468, 13'sd2172, 13'sd2735}, {12'sd-1931, 11'sd-829, 12'sd-1423}},
{{12'sd-2009, 13'sd2540, 13'sd2129}, {12'sd1361, 11'sd-870, 12'sd1344}, {10'sd386, 11'sd-739, 13'sd2409}},
{{12'sd-1213, 13'sd-2920, 12'sd1938}, {13'sd-2388, 11'sd797, 12'sd-1522}, {12'sd1427, 10'sd442, 11'sd-613}}},
{
{{13'sd2388, 12'sd1046, 12'sd1570}, {12'sd1804, 10'sd-287, 13'sd2123}, {13'sd-2273, 12'sd-1261, 13'sd2051}},
{{12'sd1297, 5'sd11, 13'sd-2252}, {12'sd-1684, 11'sd773, 12'sd1210}, {11'sd-543, 12'sd-1517, 11'sd714}},
{{12'sd1181, 12'sd-1152, 13'sd-2412}, {12'sd1069, 12'sd-1547, 9'sd-210}, {12'sd1678, 12'sd-1061, 11'sd719}},
{{13'sd-2270, 13'sd2468, 12'sd-1257}, {12'sd-1041, 11'sd-769, 13'sd2359}, {13'sd-2401, 11'sd-893, 1'sd0}},
{{11'sd947, 13'sd3229, 10'sd505}, {14'sd4921, 11'sd838, 13'sd2082}, {12'sd1520, 12'sd1869, 10'sd491}},
{{12'sd1636, 12'sd1053, 11'sd751}, {12'sd-1731, 7'sd-47, 11'sd-768}, {13'sd-2838, 12'sd-1820, 13'sd2059}},
{{10'sd-330, 13'sd3407, 13'sd2586}, {12'sd1526, 10'sd287, 12'sd1165}, {13'sd-2506, 13'sd-2399, 11'sd969}},
{{12'sd-1830, 11'sd968, 13'sd2091}, {13'sd-2347, 13'sd2532, 11'sd512}, {8'sd-101, 11'sd-716, 13'sd-2553}},
{{10'sd-509, 13'sd-2549, 13'sd-2391}, {13'sd2278, 11'sd-517, 12'sd-1101}, {11'sd-675, 11'sd558, 13'sd-2495}},
{{12'sd1779, 7'sd-50, 12'sd1081}, {10'sd-402, 11'sd-821, 13'sd-2157}, {12'sd-1042, 9'sd192, 12'sd1646}},
{{10'sd256, 10'sd-401, 12'sd-1580}, {13'sd-2089, 13'sd-2497, 12'sd-1547}, {13'sd2456, 11'sd890, 12'sd1533}},
{{12'sd1945, 12'sd-1415, 11'sd-810}, {12'sd1661, 12'sd-1909, 11'sd873}, {13'sd2138, 13'sd-2233, 11'sd643}},
{{12'sd1773, 9'sd-152, 12'sd1323}, {11'sd-938, 9'sd227, 11'sd869}, {8'sd-114, 13'sd2581, 11'sd788}},
{{7'sd45, 13'sd-2290, 9'sd247}, {11'sd924, 13'sd-2375, 12'sd-2028}, {10'sd-346, 12'sd-1260, 13'sd2149}},
{{12'sd1592, 12'sd1987, 12'sd1732}, {13'sd3775, 11'sd-829, 9'sd148}, {12'sd1841, 13'sd3179, 12'sd1504}},
{{10'sd-295, 12'sd1125, 13'sd-2754}, {12'sd1186, 2'sd1, 12'sd-1537}, {11'sd-807, 11'sd816, 13'sd2566}},
{{12'sd-1463, 13'sd-2086, 10'sd-291}, {12'sd-1209, 13'sd2072, 13'sd-2528}, {13'sd2393, 10'sd462, 11'sd627}},
{{8'sd-99, 12'sd-1288, 13'sd3028}, {8'sd-109, 12'sd-1599, 11'sd-794}, {12'sd1352, 12'sd-1394, 10'sd-464}},
{{12'sd-1498, 12'sd-1087, 11'sd598}, {11'sd-751, 11'sd933, 12'sd-1591}, {13'sd-2155, 11'sd752, 13'sd-2453}},
{{12'sd-1318, 12'sd-2042, 10'sd-468}, {13'sd-2706, 11'sd885, 13'sd2203}, {12'sd-1508, 13'sd2243, 13'sd-2431}},
{{12'sd1094, 11'sd-853, 12'sd1732}, {12'sd-1140, 12'sd1448, 12'sd1106}, {12'sd1376, 11'sd539, 13'sd-2455}},
{{11'sd-744, 11'sd738, 12'sd1361}, {12'sd-1799, 12'sd-1756, 13'sd-2190}, {12'sd1715, 11'sd-618, 13'sd-2538}},
{{10'sd-401, 12'sd-1623, 12'sd1123}, {13'sd2265, 13'sd2178, 12'sd-1958}, {12'sd-1135, 12'sd-1966, 11'sd-730}},
{{11'sd618, 12'sd2015, 7'sd49}, {13'sd-2329, 13'sd-2372, 13'sd-2096}, {13'sd-2347, 9'sd240, 12'sd-1134}},
{{13'sd-2242, 13'sd2832, 13'sd2449}, {12'sd1066, 12'sd-1466, 6'sd-29}, {12'sd-1854, 11'sd850, 11'sd534}},
{{11'sd-669, 13'sd2205, 13'sd2739}, {13'sd2761, 9'sd-207, 10'sd-382}, {12'sd-1524, 12'sd-1692, 11'sd-627}},
{{11'sd746, 9'sd-196, 12'sd1072}, {11'sd-799, 11'sd-1015, 6'sd-31}, {12'sd-1368, 11'sd-772, 13'sd-2546}},
{{13'sd2568, 12'sd1512, 13'sd2294}, {9'sd-155, 11'sd-760, 12'sd-1173}, {13'sd2522, 12'sd1211, 11'sd-537}},
{{12'sd1245, 13'sd2269, 12'sd1501}, {12'sd-1843, 13'sd-2190, 12'sd1348}, {12'sd1074, 12'sd-1100, 12'sd1716}},
{{12'sd-1039, 12'sd-1689, 13'sd2367}, {10'sd361, 13'sd-2267, 12'sd1298}, {13'sd2130, 11'sd-650, 11'sd638}},
{{13'sd2662, 13'sd2407, 13'sd2568}, {11'sd-910, 11'sd746, 11'sd-627}, {11'sd-738, 11'sd-777, 12'sd-1685}},
{{12'sd1066, 12'sd1335, 13'sd2349}, {12'sd1918, 12'sd-1385, 5'sd-14}, {12'sd1431, 13'sd-2304, 12'sd1168}},
{{13'sd2658, 12'sd1971, 12'sd-1194}, {11'sd943, 13'sd-2626, 11'sd996}, {11'sd-917, 12'sd1557, 12'sd-1873}},
{{12'sd-1904, 10'sd262, 13'sd-2806}, {11'sd-929, 12'sd-1641, 8'sd-113}, {11'sd825, 11'sd708, 12'sd2026}},
{{12'sd-1686, 12'sd-1839, 12'sd1211}, {11'sd-574, 13'sd-2086, 12'sd-2017}, {12'sd1427, 12'sd-2019, 13'sd-2980}},
{{12'sd1645, 12'sd-1746, 12'sd-1025}, {13'sd-2103, 11'sd536, 11'sd516}, {8'sd-74, 12'sd-1200, 12'sd1279}},
{{9'sd190, 9'sd-161, 14'sd-4574}, {12'sd-1674, 1'sd0, 13'sd-3187}, {12'sd1840, 13'sd-3118, 12'sd-1177}},
{{11'sd609, 13'sd2788, 11'sd725}, {12'sd1794, 11'sd601, 12'sd1460}, {13'sd2494, 12'sd-2015, 12'sd-1441}},
{{13'sd2191, 13'sd-2495, 12'sd-1897}, {7'sd-47, 13'sd2400, 13'sd-2065}, {10'sd438, 12'sd1310, 13'sd2194}},
{{11'sd865, 12'sd-1032, 13'sd-2182}, {12'sd1821, 12'sd-1658, 10'sd470}, {13'sd2688, 12'sd1159, 12'sd1106}},
{{10'sd-473, 13'sd2162, 10'sd-332}, {12'sd1227, 8'sd-85, 9'sd204}, {12'sd1716, 10'sd-337, 12'sd-1820}},
{{11'sd755, 12'sd-1838, 12'sd-1110}, {11'sd766, 11'sd871, 10'sd380}, {12'sd1734, 12'sd1314, 13'sd3654}},
{{9'sd-213, 9'sd-138, 12'sd1064}, {12'sd-1425, 12'sd1140, 12'sd1236}, {11'sd882, 13'sd-2370, 11'sd-994}},
{{12'sd-1400, 12'sd-1295, 12'sd-1338}, {12'sd1480, 13'sd2247, 12'sd1458}, {12'sd1124, 11'sd-958, 13'sd3039}},
{{12'sd1383, 13'sd2368, 12'sd1681}, {10'sd-422, 12'sd1235, 11'sd586}, {11'sd-627, 9'sd152, 12'sd-1659}},
{{10'sd-257, 8'sd-96, 11'sd-652}, {13'sd-2397, 13'sd2348, 13'sd-2513}, {11'sd725, 9'sd213, 12'sd1633}},
{{13'sd-2609, 12'sd1649, 12'sd1904}, {13'sd-2276, 8'sd95, 10'sd-391}, {10'sd384, 7'sd37, 12'sd-2044}},
{{12'sd1425, 12'sd1267, 11'sd874}, {13'sd3010, 12'sd1669, 12'sd1698}, {12'sd1640, 12'sd-1708, 13'sd2473}},
{{11'sd-802, 4'sd-4, 12'sd1269}, {13'sd2401, 11'sd-594, 12'sd-1908}, {12'sd1394, 13'sd-3145, 13'sd-2854}},
{{12'sd2004, 13'sd-3069, 13'sd-2180}, {6'sd-16, 12'sd-1972, 11'sd-814}, {12'sd1851, 13'sd-3286, 8'sd81}},
{{12'sd-1341, 13'sd-2367, 12'sd1524}, {11'sd-859, 11'sd-669, 12'sd1145}, {12'sd-1097, 10'sd286, 13'sd2363}},
{{7'sd48, 8'sd-77, 12'sd-1846}, {10'sd-317, 12'sd1325, 13'sd2342}, {11'sd-796, 13'sd2277, 10'sd281}},
{{9'sd187, 10'sd-476, 12'sd1537}, {12'sd-1851, 12'sd-1414, 13'sd-2057}, {13'sd2247, 13'sd2926, 13'sd2349}},
{{11'sd967, 12'sd-1107, 11'sd648}, {13'sd-2529, 13'sd2293, 12'sd-1267}, {12'sd-1609, 12'sd1356, 11'sd673}},
{{13'sd2898, 10'sd-437, 11'sd516}, {10'sd-467, 13'sd2717, 12'sd2039}, {7'sd-58, 9'sd-168, 9'sd-176}},
{{12'sd1844, 11'sd-538, 6'sd27}, {13'sd2119, 12'sd-1038, 12'sd1628}, {9'sd173, 10'sd354, 13'sd-3106}},
{{11'sd618, 13'sd2516, 14'sd4490}, {11'sd-789, 13'sd2129, 11'sd662}, {13'sd3975, 14'sd4684, 13'sd2332}},
{{12'sd1369, 12'sd-1907, 13'sd2200}, {12'sd-1155, 12'sd-1361, 13'sd2466}, {10'sd497, 12'sd1142, 9'sd-144}},
{{13'sd2140, 12'sd1657, 12'sd-1510}, {13'sd2447, 13'sd2679, 13'sd2948}, {13'sd-2502, 13'sd2093, 13'sd2670}},
{{11'sd-918, 10'sd-392, 13'sd2258}, {10'sd450, 12'sd1730, 10'sd293}, {11'sd960, 13'sd-2440, 11'sd-609}},
{{13'sd2217, 12'sd1338, 10'sd280}, {11'sd-867, 12'sd1889, 11'sd-585}, {12'sd-1460, 10'sd465, 12'sd1119}},
{{12'sd2047, 10'sd-375, 11'sd-931}, {12'sd1201, 12'sd-1159, 13'sd-2517}, {13'sd2160, 12'sd1267, 11'sd-829}},
{{13'sd2830, 12'sd-1218, 13'sd-2679}, {13'sd2275, 12'sd-1882, 13'sd-2299}, {13'sd2879, 13'sd-2776, 9'sd-130}},
{{12'sd1084, 12'sd1680, 10'sd-392}, {12'sd-1223, 9'sd144, 12'sd-1173}, {12'sd1683, 12'sd1228, 12'sd1245}}},
{
{{13'sd2632, 12'sd2005, 13'sd-2970}, {12'sd1099, 11'sd-972, 12'sd1588}, {12'sd-1854, 10'sd-504, 13'sd-2574}},
{{13'sd2916, 12'sd-1803, 9'sd-188}, {11'sd1007, 12'sd-1109, 9'sd251}, {11'sd-638, 12'sd1036, 11'sd-883}},
{{10'sd-262, 12'sd-1939, 12'sd1100}, {13'sd-2695, 13'sd-2143, 12'sd-1600}, {12'sd1707, 10'sd305, 12'sd-1047}},
{{11'sd518, 12'sd-1063, 12'sd1057}, {10'sd408, 12'sd1444, 12'sd-2007}, {12'sd1110, 11'sd-837, 12'sd-1499}},
{{12'sd1227, 11'sd-1001, 13'sd3093}, {13'sd3713, 10'sd-431, 10'sd-481}, {13'sd3825, 11'sd764, 12'sd1124}},
{{11'sd-681, 12'sd1252, 13'sd-2397}, {13'sd-2257, 12'sd-1125, 10'sd-443}, {12'sd1317, 12'sd1459, 11'sd-923}},
{{10'sd-445, 12'sd1058, 13'sd-3352}, {13'sd3575, 13'sd2905, 12'sd-1030}, {12'sd-2006, 11'sd-838, 10'sd-285}},
{{10'sd-382, 11'sd978, 13'sd-3246}, {8'sd125, 12'sd-1800, 12'sd-1332}, {10'sd-504, 11'sd-607, 10'sd490}},
{{12'sd1517, 11'sd-627, 12'sd1889}, {13'sd-2402, 13'sd2494, 13'sd2387}, {6'sd-17, 11'sd-845, 13'sd2399}},
{{12'sd-1085, 10'sd428, 13'sd-2363}, {13'sd-2637, 12'sd1717, 12'sd1411}, {12'sd-1091, 12'sd-1194, 13'sd-2729}},
{{13'sd-2854, 11'sd601, 12'sd-1640}, {10'sd-478, 10'sd361, 12'sd1027}, {12'sd-1498, 11'sd723, 12'sd-1713}},
{{13'sd-2454, 13'sd2131, 12'sd1529}, {11'sd701, 12'sd-1521, 13'sd-2541}, {12'sd-1173, 13'sd-2320, 11'sd-612}},
{{12'sd1100, 11'sd-941, 11'sd-512}, {12'sd-1529, 13'sd2420, 12'sd-2030}, {9'sd-137, 12'sd-1207, 12'sd-1899}},
{{11'sd985, 11'sd800, 12'sd1414}, {11'sd-793, 12'sd-1925, 12'sd-1587}, {12'sd1081, 13'sd2258, 9'sd137}},
{{12'sd1958, 7'sd-60, 13'sd3000}, {11'sd-837, 13'sd3539, 13'sd2717}, {11'sd-838, 12'sd1194, 14'sd5111}},
{{12'sd1523, 12'sd-1694, 8'sd86}, {11'sd557, 12'sd1333, 12'sd1572}, {12'sd1262, 11'sd770, 12'sd-1976}},
{{10'sd290, 11'sd-933, 11'sd577}, {11'sd579, 12'sd1210, 10'sd-406}, {13'sd2717, 10'sd356, 9'sd164}},
{{9'sd-198, 12'sd1226, 9'sd-190}, {10'sd301, 13'sd2662, 10'sd-322}, {13'sd2713, 10'sd-457, 13'sd2971}},
{{11'sd-951, 13'sd-2429, 8'sd105}, {12'sd-1854, 13'sd2074, 9'sd242}, {12'sd1611, 12'sd1200, 11'sd711}},
{{12'sd1086, 12'sd-1730, 10'sd335}, {9'sd-254, 10'sd-401, 13'sd-2497}, {8'sd-101, 9'sd230, 11'sd-805}},
{{13'sd-2352, 12'sd1939, 12'sd1834}, {9'sd203, 13'sd2057, 13'sd2129}, {13'sd-2560, 7'sd-39, 12'sd-1529}},
{{13'sd-2661, 12'sd-1052, 10'sd-376}, {12'sd1586, 13'sd2613, 13'sd-2136}, {12'sd1439, 7'sd-42, 13'sd-2477}},
{{12'sd-1486, 7'sd-40, 13'sd2387}, {12'sd-2032, 13'sd-2302, 9'sd227}, {13'sd2142, 12'sd-1088, 12'sd-1337}},
{{12'sd-1716, 9'sd-151, 11'sd780}, {13'sd2570, 11'sd585, 13'sd2105}, {13'sd-2412, 13'sd2425, 12'sd-1345}},
{{10'sd-453, 12'sd1132, 12'sd-1673}, {13'sd-2109, 10'sd-368, 11'sd574}, {13'sd2506, 10'sd430, 9'sd169}},
{{11'sd808, 13'sd2870, 11'sd-957}, {9'sd226, 13'sd-2246, 10'sd410}, {13'sd2260, 10'sd352, 12'sd1324}},
{{13'sd-2324, 8'sd-102, 11'sd-754}, {12'sd-1571, 9'sd-203, 13'sd-2598}, {13'sd-3020, 11'sd-670, 11'sd-894}},
{{13'sd2244, 13'sd3144, 13'sd3477}, {10'sd373, 10'sd-298, 12'sd-1889}, {12'sd-1563, 9'sd220, 13'sd2135}},
{{10'sd471, 11'sd619, 12'sd-1359}, {11'sd911, 7'sd45, 9'sd-136}, {12'sd-1233, 12'sd1855, 13'sd2148}},
{{12'sd-1211, 12'sd-1306, 9'sd201}, {9'sd-230, 13'sd2213, 13'sd-2357}, {12'sd-1574, 13'sd-2342, 10'sd-408}},
{{8'sd-116, 8'sd76, 12'sd-1400}, {13'sd2128, 11'sd825, 13'sd2269}, {9'sd-245, 13'sd2108, 9'sd244}},
{{12'sd1224, 13'sd2099, 13'sd2714}, {11'sd-513, 9'sd-204, 12'sd1075}, {13'sd-2150, 10'sd350, 13'sd2426}},
{{9'sd255, 13'sd2054, 10'sd-295}, {12'sd-1759, 11'sd992, 13'sd-2105}, {9'sd-223, 12'sd-1311, 7'sd43}},
{{12'sd1032, 12'sd-1105, 13'sd2552}, {12'sd1623, 13'sd2510, 13'sd3151}, {12'sd1665, 12'sd-1061, 12'sd1802}},
{{12'sd1790, 13'sd-2396, 9'sd-237}, {10'sd-410, 10'sd295, 13'sd2205}, {12'sd1249, 12'sd-1676, 13'sd2236}},
{{12'sd-1351, 11'sd855, 8'sd68}, {13'sd-2188, 10'sd-463, 10'sd-482}, {11'sd-674, 12'sd-1241, 12'sd1554}},
{{11'sd-873, 8'sd-73, 13'sd-2339}, {12'sd1896, 9'sd214, 13'sd-2076}, {12'sd1994, 13'sd-3324, 11'sd945}},
{{12'sd1722, 12'sd1443, 7'sd61}, {12'sd-1996, 9'sd129, 11'sd-675}, {12'sd-1978, 13'sd2722, 11'sd740}},
{{9'sd245, 12'sd-1690, 12'sd1880}, {12'sd1988, 11'sd-649, 11'sd-830}, {13'sd-2696, 11'sd650, 9'sd245}},
{{13'sd2262, 12'sd1124, 13'sd2611}, {13'sd-2733, 11'sd749, 12'sd-2027}, {11'sd570, 13'sd2304, 11'sd-925}},
{{8'sd101, 12'sd-1757, 12'sd-1061}, {11'sd-841, 10'sd-381, 12'sd-1979}, {12'sd1597, 12'sd-1886, 12'sd-1974}},
{{8'sd-88, 12'sd-1158, 12'sd1717}, {12'sd1126, 12'sd-1504, 12'sd-1699}, {11'sd1013, 12'sd-1107, 13'sd2087}},
{{12'sd-1453, 13'sd2981, 12'sd1803}, {11'sd558, 12'sd-1427, 12'sd1763}, {13'sd-3401, 11'sd-939, 13'sd3021}},
{{8'sd109, 9'sd208, 13'sd-2507}, {11'sd559, 13'sd2977, 13'sd-3459}, {10'sd-289, 10'sd472, 12'sd1193}},
{{13'sd-2329, 13'sd-2133, 10'sd370}, {10'sd-509, 12'sd1205, 10'sd259}, {12'sd-1052, 13'sd-2812, 12'sd-1499}},
{{11'sd589, 11'sd872, 10'sd-353}, {9'sd140, 12'sd1929, 9'sd200}, {10'sd-443, 13'sd-2177, 10'sd-461}},
{{10'sd373, 11'sd-661, 12'sd-1927}, {10'sd294, 13'sd-2921, 13'sd2177}, {12'sd1167, 12'sd1956, 13'sd2500}},
{{12'sd1406, 13'sd2569, 13'sd2192}, {12'sd1039, 10'sd332, 13'sd3057}, {9'sd-182, 9'sd224, 11'sd-547}},
{{12'sd1326, 11'sd895, 13'sd-2346}, {7'sd-61, 10'sd276, 13'sd2121}, {12'sd-1851, 11'sd889, 13'sd-2596}},
{{11'sd-598, 12'sd-1884, 11'sd-1017}, {13'sd-3206, 11'sd776, 11'sd781}, {13'sd2934, 10'sd-451, 12'sd1382}},
{{10'sd275, 13'sd-2062, 9'sd236}, {11'sd-588, 10'sd-340, 12'sd-1733}, {12'sd1480, 11'sd736, 12'sd1122}},
{{11'sd-979, 12'sd-1417, 12'sd-1497}, {13'sd-2154, 9'sd131, 13'sd-2259}, {11'sd-685, 11'sd565, 11'sd-578}},
{{11'sd-669, 10'sd325, 12'sd-1811}, {7'sd57, 12'sd-1649, 13'sd2775}, {12'sd1729, 13'sd2572, 12'sd-1986}},
{{10'sd383, 12'sd-1463, 10'sd-406}, {11'sd-709, 11'sd887, 13'sd2534}, {10'sd-456, 13'sd2188, 11'sd-592}},
{{13'sd2436, 12'sd-1539, 13'sd2165}, {9'sd203, 12'sd-1490, 12'sd1990}, {11'sd1012, 10'sd326, 12'sd1645}},
{{11'sd-748, 5'sd9, 13'sd-2242}, {12'sd1125, 11'sd-557, 13'sd-2622}, {12'sd1819, 12'sd2012, 12'sd1858}},
{{12'sd1325, 10'sd-271, 13'sd-2309}, {13'sd2231, 8'sd-83, 7'sd-61}, {13'sd3116, 13'sd-2341, 13'sd-2338}},
{{11'sd-847, 11'sd771, 10'sd-349}, {13'sd2358, 11'sd-969, 12'sd-1415}, {12'sd-1629, 11'sd551, 11'sd801}},
{{12'sd1233, 12'sd1175, 12'sd1869}, {11'sd657, 13'sd2268, 11'sd596}, {11'sd853, 12'sd1246, 11'sd547}},
{{11'sd-781, 13'sd3035, 14'sd4186}, {12'sd1640, 9'sd-165, 13'sd2118}, {11'sd626, 12'sd-1622, 12'sd2006}},
{{11'sd893, 13'sd2385, 9'sd180}, {10'sd508, 12'sd-1931, 12'sd1589}, {9'sd236, 11'sd741, 11'sd-922}},
{{13'sd2267, 9'sd176, 10'sd-271}, {12'sd-1599, 12'sd-1640, 12'sd-1471}, {8'sd115, 13'sd-2396, 11'sd879}},
{{12'sd-1678, 12'sd1139, 13'sd-2770}, {12'sd-1906, 9'sd-240, 13'sd-2628}, {9'sd244, 11'sd-986, 10'sd433}},
{{10'sd-337, 12'sd-1183, 6'sd19}, {9'sd-232, 13'sd2309, 7'sd34}, {11'sd838, 13'sd2073, 12'sd1708}}},
{
{{12'sd1601, 12'sd-1293, 12'sd-1149}, {11'sd753, 12'sd-1233, 11'sd540}, {12'sd-1175, 11'sd-797, 11'sd899}},
{{13'sd2449, 12'sd1216, 12'sd-1257}, {13'sd2082, 13'sd2262, 13'sd2566}, {12'sd1675, 13'sd2124, 12'sd1775}},
{{11'sd686, 13'sd2850, 12'sd-1450}, {10'sd450, 11'sd-628, 12'sd1352}, {11'sd576, 12'sd-1106, 12'sd1653}},
{{13'sd2136, 11'sd-668, 13'sd2260}, {13'sd-2917, 13'sd-3093, 13'sd-2988}, {11'sd564, 12'sd-1313, 11'sd-803}},
{{13'sd3484, 14'sd4199, 12'sd1668}, {13'sd-2882, 12'sd-1251, 10'sd-406}, {12'sd-1864, 8'sd82, 11'sd-924}},
{{13'sd2622, 12'sd1083, 13'sd2412}, {11'sd-607, 12'sd1463, 10'sd311}, {13'sd2944, 11'sd840, 12'sd-1724}},
{{10'sd-324, 12'sd1603, 11'sd553}, {13'sd-2742, 11'sd843, 13'sd-2378}, {12'sd1412, 12'sd-1454, 14'sd-4180}},
{{9'sd234, 13'sd-2471, 12'sd1598}, {12'sd-2047, 11'sd-535, 11'sd-513}, {8'sd-104, 13'sd2440, 9'sd-242}},
{{12'sd-1930, 12'sd-1781, 12'sd-1460}, {10'sd290, 8'sd76, 13'sd2373}, {12'sd1083, 12'sd1473, 11'sd-576}},
{{12'sd1579, 13'sd-2218, 12'sd-1419}, {11'sd665, 13'sd-2911, 12'sd1694}, {11'sd-826, 6'sd-26, 9'sd-148}},
{{10'sd-339, 12'sd-1780, 12'sd1396}, {8'sd-91, 12'sd1568, 10'sd502}, {10'sd324, 12'sd-2002, 9'sd144}},
{{10'sd-474, 11'sd-748, 12'sd-1519}, {11'sd673, 11'sd582, 9'sd198}, {12'sd1992, 11'sd-554, 8'sd124}},
{{12'sd-1289, 10'sd-340, 11'sd828}, {11'sd-913, 13'sd-2054, 11'sd540}, {10'sd-327, 13'sd-3997, 11'sd-895}},
{{13'sd-2760, 13'sd2521, 13'sd2614}, {13'sd-2460, 12'sd1437, 12'sd1459}, {13'sd2293, 13'sd-2306, 13'sd2896}},
{{11'sd691, 12'sd-1621, 13'sd-2805}, {9'sd224, 12'sd1881, 13'sd-3290}, {11'sd-643, 12'sd-1067, 10'sd494}},
{{12'sd-1678, 12'sd1985, 13'sd-2152}, {12'sd2023, 13'sd2963, 12'sd-1660}, {13'sd2459, 12'sd-1921, 12'sd1667}},
{{12'sd-1334, 12'sd1576, 12'sd1209}, {9'sd230, 13'sd-2820, 11'sd894}, {13'sd2535, 12'sd1505, 12'sd1102}},
{{12'sd1048, 8'sd114, 11'sd-580}, {11'sd-908, 13'sd2378, 11'sd639}, {13'sd-2329, 12'sd-1262, 9'sd-163}},
{{11'sd939, 13'sd2432, 10'sd-457}, {11'sd-867, 12'sd-1087, 12'sd1346}, {12'sd2009, 12'sd1224, 13'sd-2466}},
{{13'sd-2090, 13'sd-2135, 10'sd258}, {12'sd1667, 12'sd1087, 11'sd662}, {11'sd-939, 12'sd1990, 7'sd-41}},
{{8'sd79, 13'sd2381, 13'sd-3009}, {12'sd1873, 12'sd-1741, 8'sd-113}, {12'sd-1233, 11'sd-982, 12'sd-1397}},
{{9'sd-193, 8'sd66, 13'sd2522}, {10'sd426, 10'sd-447, 11'sd1017}, {11'sd639, 12'sd-1314, 10'sd-398}},
{{13'sd-2692, 12'sd1100, 13'sd2239}, {12'sd1878, 11'sd-900, 11'sd945}, {7'sd-59, 10'sd287, 10'sd-362}},
{{11'sd564, 13'sd2062, 11'sd-960}, {12'sd-1159, 13'sd2162, 11'sd660}, {12'sd-1643, 8'sd73, 12'sd1258}},
{{11'sd580, 13'sd-2409, 12'sd-1187}, {12'sd-1907, 9'sd162, 11'sd-516}, {11'sd860, 11'sd-561, 11'sd542}},
{{12'sd-1086, 12'sd1817, 13'sd2610}, {13'sd2170, 9'sd222, 12'sd1372}, {12'sd-1197, 12'sd-2024, 11'sd659}},
{{13'sd3487, 6'sd30, 11'sd868}, {3'sd-2, 9'sd151, 10'sd-423}, {13'sd2876, 12'sd1377, 12'sd-1146}},
{{12'sd1923, 12'sd1709, 12'sd2043}, {10'sd484, 12'sd-1519, 12'sd1956}, {12'sd-1761, 13'sd-3572, 10'sd-330}},
{{9'sd242, 12'sd1747, 12'sd-1572}, {11'sd-573, 12'sd-1625, 12'sd1776}, {12'sd-1953, 13'sd2388, 11'sd721}},
{{13'sd2406, 12'sd-1045, 13'sd-2426}, {10'sd-442, 12'sd-1252, 12'sd-1672}, {12'sd1630, 12'sd-1307, 13'sd2924}},
{{10'sd-280, 7'sd-59, 12'sd1653}, {12'sd-1857, 12'sd-1741, 12'sd1207}, {13'sd2124, 12'sd1969, 12'sd-1503}},
{{13'sd2121, 12'sd1412, 12'sd1558}, {11'sd802, 7'sd40, 12'sd1874}, {11'sd-988, 9'sd-225, 8'sd72}},
{{9'sd212, 12'sd-1235, 11'sd520}, {12'sd1829, 12'sd-1675, 12'sd1706}, {12'sd-1924, 7'sd60, 13'sd2729}},
{{13'sd2693, 12'sd-1107, 9'sd-159}, {10'sd-330, 12'sd1643, 10'sd-507}, {9'sd146, 12'sd-1209, 13'sd2434}},
{{13'sd2243, 12'sd-1720, 12'sd1763}, {13'sd2766, 13'sd3245, 12'sd1524}, {13'sd3248, 11'sd895, 13'sd3759}},
{{11'sd-921, 12'sd1732, 12'sd2007}, {13'sd2186, 13'sd2079, 11'sd-1003}, {13'sd2476, 13'sd2107, 10'sd422}},
{{13'sd2818, 12'sd-1572, 13'sd-3332}, {13'sd3292, 10'sd363, 10'sd-442}, {12'sd2033, 10'sd373, 13'sd3322}},
{{13'sd2935, 12'sd1372, 12'sd1793}, {12'sd1265, 10'sd324, 5'sd11}, {11'sd-907, 13'sd2069, 10'sd-488}},
{{9'sd169, 11'sd956, 13'sd2815}, {10'sd492, 11'sd1008, 13'sd-2388}, {11'sd1015, 11'sd988, 13'sd-2931}},
{{12'sd1801, 12'sd1104, 11'sd895}, {12'sd-1945, 12'sd1174, 13'sd2155}, {13'sd-2055, 11'sd-694, 12'sd-1858}},
{{13'sd2837, 12'sd-1991, 9'sd-160}, {13'sd2530, 8'sd83, 12'sd-1517}, {11'sd700, 11'sd531, 12'sd1678}},
{{13'sd2338, 12'sd-1592, 12'sd1625}, {11'sd1023, 12'sd-1418, 13'sd2338}, {10'sd399, 11'sd694, 13'sd-2446}},
{{12'sd1309, 10'sd301, 12'sd1991}, {11'sd887, 12'sd-1990, 10'sd509}, {12'sd-1610, 10'sd468, 12'sd1250}},
{{13'sd3601, 13'sd3325, 12'sd1460}, {12'sd1974, 12'sd1401, 12'sd-1493}, {10'sd487, 11'sd622, 12'sd-1591}},
{{12'sd1129, 13'sd-2566, 11'sd985}, {13'sd2749, 12'sd1150, 12'sd1725}, {13'sd2434, 13'sd-2288, 12'sd-1215}},
{{11'sd731, 12'sd-1400, 12'sd-1387}, {13'sd2427, 13'sd2508, 12'sd-1352}, {11'sd-568, 12'sd1213, 12'sd1125}},
{{10'sd360, 12'sd-1461, 11'sd-993}, {13'sd2357, 11'sd909, 13'sd3077}, {9'sd158, 1'sd0, 13'sd2111}},
{{12'sd1556, 10'sd-334, 10'sd345}, {10'sd-367, 12'sd-1173, 10'sd-276}, {11'sd-761, 12'sd-1287, 13'sd2644}},
{{11'sd877, 13'sd2746, 13'sd-2569}, {13'sd3747, 11'sd-618, 13'sd-2883}, {13'sd3489, 12'sd-1200, 8'sd113}},
{{12'sd-1683, 13'sd-3028, 12'sd-1899}, {10'sd417, 7'sd42, 11'sd-653}, {12'sd-1898, 11'sd850, 11'sd1009}},
{{13'sd2173, 13'sd2741, 13'sd2455}, {8'sd-76, 12'sd-1833, 13'sd2409}, {9'sd-205, 13'sd2070, 13'sd2440}},
{{10'sd-294, 13'sd-2656, 11'sd813}, {11'sd-851, 12'sd-1538, 10'sd-502}, {12'sd-1617, 12'sd1291, 13'sd-3225}},
{{11'sd745, 13'sd-2467, 12'sd1363}, {13'sd-2396, 9'sd-177, 12'sd-1596}, {12'sd-1514, 13'sd-2929, 11'sd-938}},
{{13'sd2226, 13'sd2313, 11'sd982}, {11'sd-955, 12'sd-1637, 11'sd-863}, {13'sd3367, 12'sd-1256, 12'sd-1635}},
{{12'sd-1385, 11'sd881, 13'sd2579}, {10'sd-309, 8'sd-114, 11'sd922}, {11'sd928, 8'sd-91, 9'sd235}},
{{11'sd514, 10'sd-388, 13'sd-2219}, {12'sd1370, 10'sd297, 12'sd1140}, {11'sd-704, 12'sd-1837, 13'sd-2462}},
{{12'sd-1554, 13'sd2207, 8'sd-110}, {13'sd-3789, 12'sd-1760, 13'sd-2791}, {13'sd-3716, 13'sd-3927, 13'sd-3120}},
{{13'sd2556, 11'sd992, 13'sd2299}, {13'sd2309, 13'sd2200, 10'sd366}, {11'sd590, 9'sd158, 11'sd963}},
{{12'sd1361, 11'sd830, 11'sd-732}, {13'sd3068, 11'sd998, 11'sd665}, {5'sd-12, 12'sd-1363, 9'sd-214}},
{{13'sd2894, 12'sd1958, 12'sd-1313}, {13'sd3854, 13'sd3111, 12'sd-1950}, {13'sd3620, 10'sd-335, 12'sd1514}},
{{11'sd519, 13'sd2334, 6'sd18}, {13'sd-2486, 12'sd-1138, 10'sd-361}, {12'sd1085, 12'sd1879, 13'sd-2147}},
{{8'sd-68, 12'sd-1893, 13'sd-2459}, {12'sd-1572, 10'sd459, 13'sd-2187}, {12'sd-1538, 10'sd-322, 13'sd-3358}},
{{12'sd-1296, 12'sd-1233, 12'sd-1832}, {12'sd-1443, 11'sd-777, 13'sd2084}, {12'sd1119, 12'sd-1733, 13'sd2472}},
{{12'sd-1415, 13'sd-2177, 12'sd-1162}, {12'sd1974, 13'sd-2712, 12'sd-1707}, {12'sd1102, 12'sd1136, 13'sd-3015}}},
{
{{13'sd-2162, 11'sd-615, 11'sd-618}, {8'sd-88, 13'sd-2524, 11'sd861}, {13'sd-2521, 12'sd1398, 13'sd-2808}},
{{12'sd1924, 12'sd1879, 11'sd515}, {13'sd-2076, 12'sd1904, 11'sd-766}, {12'sd-1046, 12'sd1965, 6'sd18}},
{{13'sd-2547, 11'sd-791, 12'sd1412}, {13'sd2170, 13'sd2538, 10'sd-433}, {9'sd171, 10'sd327, 13'sd-2295}},
{{12'sd-1037, 10'sd306, 5'sd-11}, {10'sd-413, 11'sd632, 12'sd1224}, {13'sd2482, 13'sd-2393, 11'sd-951}},
{{12'sd-1446, 12'sd1688, 11'sd886}, {13'sd-3923, 8'sd-94, 10'sd333}, {11'sd545, 2'sd-1, 13'sd-2289}},
{{10'sd-354, 11'sd-908, 13'sd-2771}, {12'sd1799, 13'sd-2292, 11'sd-895}, {12'sd1788, 11'sd-920, 13'sd2199}},
{{13'sd2145, 10'sd-319, 8'sd112}, {6'sd28, 13'sd3446, 12'sd-1209}, {12'sd1296, 11'sd-744, 13'sd3876}},
{{11'sd-891, 10'sd-468, 13'sd-2279}, {12'sd1687, 12'sd-1417, 12'sd1047}, {12'sd1181, 13'sd2973, 12'sd-1771}},
{{11'sd-544, 11'sd-809, 12'sd-1078}, {10'sd-300, 11'sd735, 12'sd-1778}, {12'sd1802, 10'sd-471, 12'sd2005}},
{{11'sd646, 12'sd-1702, 12'sd-1584}, {13'sd-2993, 10'sd-292, 13'sd-2846}, {6'sd28, 12'sd1074, 13'sd2238}},
{{10'sd-375, 13'sd2614, 12'sd2005}, {10'sd-327, 11'sd-985, 12'sd1673}, {11'sd-758, 13'sd2368, 13'sd-2128}},
{{11'sd-539, 12'sd-1869, 8'sd84}, {13'sd-2245, 11'sd-976, 12'sd-1806}, {11'sd-652, 13'sd2292, 11'sd-702}},
{{10'sd-266, 11'sd852, 13'sd2351}, {12'sd1792, 10'sd-272, 13'sd2265}, {9'sd-248, 13'sd2124, 11'sd-689}},
{{12'sd-1625, 13'sd-2148, 13'sd2194}, {13'sd-2116, 10'sd412, 11'sd587}, {11'sd879, 12'sd1194, 13'sd2625}},
{{11'sd673, 12'sd-1884, 12'sd-1066}, {14'sd-4368, 13'sd-3226, 13'sd-2523}, {14'sd-5548, 11'sd813, 10'sd-394}},
{{13'sd2236, 12'sd-1218, 12'sd1186}, {9'sd189, 13'sd2788, 9'sd182}, {10'sd329, 12'sd-1638, 9'sd-231}},
{{10'sd-361, 10'sd411, 12'sd1756}, {13'sd2176, 13'sd2415, 12'sd-1986}, {6'sd31, 13'sd2527, 11'sd512}},
{{12'sd1245, 12'sd-1974, 13'sd2113}, {10'sd441, 10'sd-267, 12'sd-1677}, {12'sd1169, 12'sd1196, 13'sd2959}},
{{13'sd2464, 12'sd-1759, 12'sd1532}, {12'sd1407, 11'sd941, 12'sd-1432}, {12'sd1876, 10'sd-336, 12'sd1693}},
{{12'sd-1996, 12'sd1411, 12'sd-1507}, {12'sd1554, 11'sd-941, 8'sd110}, {13'sd2622, 13'sd2216, 12'sd-1623}},
{{12'sd-1345, 11'sd-786, 13'sd-2054}, {10'sd356, 12'sd-1276, 12'sd-1981}, {12'sd-1743, 11'sd-904, 7'sd-37}},
{{10'sd306, 13'sd-2605, 13'sd-2099}, {12'sd-1919, 12'sd1777, 13'sd-2542}, {13'sd2848, 11'sd514, 10'sd508}},
{{13'sd-2815, 12'sd-1467, 12'sd1042}, {12'sd1642, 12'sd1213, 12'sd1123}, {10'sd376, 10'sd-359, 13'sd2952}},
{{13'sd2535, 13'sd-2137, 11'sd933}, {12'sd1357, 12'sd-1690, 13'sd2427}, {11'sd-834, 12'sd1534, 12'sd-2007}},
{{8'sd110, 13'sd2095, 13'sd-2055}, {11'sd923, 12'sd-1066, 13'sd2982}, {11'sd718, 12'sd1879, 13'sd2324}},
{{12'sd1027, 12'sd-1801, 12'sd-1721}, {13'sd2378, 13'sd2530, 12'sd1559}, {12'sd1078, 8'sd-95, 10'sd291}},
{{14'sd4817, 13'sd3432, 12'sd1738}, {14'sd7036, 13'sd2137, 14'sd4468}, {13'sd2426, 14'sd5411, 13'sd3172}},
{{11'sd-757, 11'sd989, 11'sd-1006}, {12'sd1508, 12'sd-1963, 13'sd-2741}, {8'sd125, 11'sd-851, 11'sd-812}},
{{11'sd-979, 11'sd673, 12'sd1454}, {13'sd-2120, 10'sd-446, 12'sd-2019}, {12'sd-1957, 12'sd1406, 13'sd2300}},
{{12'sd1306, 12'sd1849, 10'sd366}, {12'sd1471, 11'sd857, 12'sd-1517}, {13'sd2067, 13'sd2431, 11'sd947}},
{{11'sd-777, 11'sd-607, 12'sd-1865}, {13'sd-2254, 10'sd-386, 9'sd-195}, {13'sd-2310, 10'sd-502, 8'sd-80}},
{{13'sd2366, 12'sd-1062, 11'sd568}, {13'sd2264, 12'sd-1450, 12'sd-1710}, {12'sd1321, 10'sd457, 12'sd1831}},
{{10'sd-313, 11'sd608, 9'sd237}, {13'sd-2269, 13'sd-2348, 11'sd-589}, {13'sd2085, 13'sd2497, 9'sd244}},
{{13'sd-2699, 12'sd-1237, 12'sd2030}, {12'sd1346, 12'sd-1873, 11'sd-923}, {12'sd-1937, 12'sd-1376, 11'sd-880}},
{{10'sd-463, 12'sd-1219, 13'sd-2110}, {13'sd-2638, 9'sd215, 12'sd-1925}, {12'sd-1308, 12'sd1138, 12'sd2026}},
{{13'sd2382, 13'sd2658, 12'sd1932}, {11'sd922, 12'sd1256, 11'sd830}, {12'sd1361, 11'sd579, 10'sd-342}},
{{13'sd3275, 8'sd-68, 9'sd160}, {11'sd731, 12'sd-1598, 12'sd1754}, {13'sd2470, 10'sd-502, 12'sd1046}},
{{13'sd2164, 11'sd-720, 13'sd-2542}, {12'sd-1504, 13'sd-2211, 11'sd861}, {13'sd-2174, 13'sd2490, 12'sd-1257}},
{{11'sd-1023, 13'sd-2311, 13'sd2886}, {13'sd2146, 12'sd1069, 8'sd-71}, {12'sd-1282, 13'sd2103, 11'sd609}},
{{10'sd-345, 11'sd-520, 11'sd896}, {10'sd483, 9'sd-193, 12'sd1782}, {13'sd-2543, 12'sd-1485, 13'sd-2220}},
{{13'sd-2086, 11'sd864, 12'sd1675}, {12'sd-1955, 9'sd-174, 11'sd696}, {13'sd2104, 8'sd100, 10'sd-348}},
{{11'sd657, 13'sd-2476, 13'sd-2722}, {12'sd1266, 12'sd1936, 12'sd1244}, {13'sd-2363, 12'sd2007, 12'sd1736}},
{{13'sd-2613, 13'sd2559, 13'sd2178}, {12'sd1107, 11'sd-958, 12'sd1750}, {12'sd-1512, 13'sd2629, 12'sd1107}},
{{13'sd3878, 13'sd3195, 13'sd-2848}, {14'sd4504, 14'sd4371, 11'sd773}, {14'sd4758, 12'sd1732, 12'sd1469}},
{{9'sd129, 13'sd2119, 13'sd-2416}, {13'sd2184, 11'sd-864, 12'sd-1863}, {12'sd1219, 12'sd1733, 12'sd1229}},
{{12'sd-1680, 13'sd-2278, 12'sd-1384}, {11'sd930, 12'sd1802, 11'sd914}, {8'sd-76, 12'sd-1807, 12'sd-1509}},
{{10'sd-277, 10'sd-375, 11'sd-997}, {10'sd-401, 13'sd-2364, 10'sd-502}, {10'sd382, 11'sd804, 10'sd-322}},
{{13'sd2917, 12'sd-1411, 13'sd-2637}, {8'sd88, 12'sd-1877, 12'sd-1722}, {12'sd-1273, 12'sd-1687, 13'sd2432}},
{{11'sd896, 10'sd-276, 12'sd-1096}, {11'sd-542, 4'sd4, 12'sd1989}, {10'sd-437, 10'sd277, 12'sd-2038}},
{{13'sd-3277, 13'sd2089, 10'sd-420}, {12'sd-1029, 13'sd-3680, 12'sd1591}, {10'sd-459, 10'sd-433, 13'sd-3256}},
{{13'sd-2488, 12'sd1224, 12'sd-1981}, {12'sd1698, 12'sd-1238, 10'sd-264}, {11'sd-993, 12'sd1168, 11'sd998}},
{{11'sd639, 13'sd2296, 12'sd1075}, {13'sd2377, 13'sd-2862, 13'sd2048}, {11'sd-513, 9'sd159, 12'sd-1469}},
{{13'sd-3611, 13'sd-2095, 8'sd122}, {12'sd1267, 10'sd464, 13'sd2292}, {13'sd-3069, 9'sd176, 13'sd-2294}},
{{4'sd-5, 9'sd-191, 11'sd-560}, {13'sd2801, 11'sd854, 13'sd2516}, {9'sd-243, 11'sd706, 12'sd1676}},
{{12'sd1717, 13'sd3244, 12'sd2017}, {12'sd-1736, 12'sd-1517, 11'sd-971}, {10'sd-429, 12'sd-1563, 8'sd80}},
{{11'sd771, 9'sd-142, 12'sd-1453}, {12'sd-2023, 12'sd1794, 12'sd1352}, {12'sd-1612, 10'sd354, 11'sd-945}},
{{12'sd1859, 10'sd-269, 12'sd1966}, {11'sd-589, 12'sd-1610, 9'sd-164}, {13'sd-3584, 13'sd-2738, 11'sd899}},
{{13'sd2593, 13'sd-2715, 11'sd557}, {13'sd-2091, 9'sd-134, 10'sd345}, {12'sd1371, 12'sd-1918, 12'sd-1307}},
{{10'sd-272, 12'sd-1516, 12'sd-1273}, {12'sd-1899, 11'sd665, 13'sd-2210}, {12'sd1740, 12'sd1794, 12'sd1613}},
{{10'sd343, 12'sd-1443, 12'sd-1391}, {12'sd1199, 11'sd-838, 13'sd2610}, {12'sd1174, 12'sd1806, 13'sd3060}},
{{12'sd-1916, 9'sd193, 12'sd-1476}, {13'sd2355, 12'sd-1156, 13'sd2795}, {12'sd1635, 12'sd-1575, 13'sd2802}},
{{13'sd-2672, 12'sd-1293, 13'sd2265}, {11'sd823, 10'sd-380, 12'sd1590}, {13'sd-2086, 13'sd-2274, 12'sd-1315}},
{{11'sd-717, 11'sd-607, 13'sd-2285}, {11'sd-1010, 9'sd-140, 8'sd-82}, {12'sd1805, 12'sd2040, 13'sd-2241}},
{{12'sd-1819, 11'sd-982, 13'sd-3060}, {11'sd921, 13'sd2053, 12'sd-1154}, {13'sd2320, 12'sd-1079, 13'sd2538}}},
{
{{11'sd716, 13'sd-2223, 12'sd1614}, {7'sd-61, 13'sd-2171, 12'sd-1289}, {11'sd-521, 13'sd-2902, 12'sd1212}},
{{11'sd-519, 11'sd706, 11'sd-649}, {13'sd2531, 12'sd1412, 12'sd1985}, {11'sd-811, 12'sd1030, 13'sd-2179}},
{{9'sd186, 8'sd-74, 12'sd1507}, {10'sd-495, 12'sd1094, 11'sd-952}, {11'sd649, 13'sd-2540, 13'sd2184}},
{{8'sd-123, 12'sd1079, 12'sd1874}, {11'sd862, 12'sd-1759, 10'sd504}, {12'sd1553, 11'sd-698, 12'sd1569}},
{{12'sd-1395, 14'sd-4172, 14'sd-4345}, {13'sd-2437, 13'sd-3154, 13'sd-3245}, {11'sd-710, 12'sd-1127, 11'sd533}},
{{12'sd-1267, 13'sd-3033, 13'sd2154}, {7'sd-32, 12'sd-1340, 12'sd1452}, {6'sd-20, 13'sd-4044, 12'sd-1632}},
{{10'sd-471, 11'sd-1012, 12'sd1143}, {13'sd-2440, 11'sd-872, 11'sd-734}, {11'sd734, 12'sd1598, 12'sd-1228}},
{{13'sd-2797, 10'sd358, 12'sd-1357}, {10'sd303, 6'sd-16, 11'sd-682}, {12'sd1527, 13'sd2434, 12'sd1083}},
{{11'sd-516, 13'sd2162, 13'sd2292}, {10'sd499, 13'sd-2214, 13'sd2281}, {13'sd-2310, 12'sd1326, 11'sd-878}},
{{12'sd1918, 12'sd1345, 13'sd-2513}, {12'sd-1819, 12'sd-1058, 13'sd-3642}, {12'sd1094, 12'sd1984, 13'sd-2984}},
{{12'sd1373, 10'sd336, 11'sd-951}, {12'sd-1781, 11'sd-813, 11'sd999}, {12'sd1815, 13'sd-2215, 10'sd-364}},
{{10'sd377, 12'sd-1182, 13'sd-2519}, {12'sd-1045, 11'sd-541, 10'sd499}, {11'sd-999, 11'sd-586, 12'sd-1683}},
{{12'sd-1419, 13'sd2511, 13'sd2609}, {10'sd-279, 11'sd-782, 12'sd1210}, {13'sd-3280, 11'sd-724, 13'sd-2110}},
{{12'sd-1692, 13'sd-3098, 12'sd-1957}, {11'sd923, 13'sd-2318, 13'sd2218}, {10'sd-464, 13'sd2054, 12'sd-1966}},
{{9'sd141, 12'sd1741, 12'sd-1581}, {13'sd2770, 4'sd-7, 12'sd-1696}, {12'sd-1714, 12'sd-1301, 11'sd647}},
{{11'sd-962, 12'sd1596, 12'sd1237}, {12'sd-1659, 12'sd-1027, 12'sd1781}, {12'sd1228, 11'sd-735, 11'sd895}},
{{13'sd-2184, 11'sd728, 11'sd-678}, {13'sd2087, 13'sd2875, 13'sd2168}, {12'sd-1967, 9'sd194, 12'sd1738}},
{{12'sd-1201, 12'sd1841, 12'sd-1127}, {13'sd-2079, 10'sd-298, 10'sd-507}, {12'sd1609, 12'sd-1852, 11'sd-610}},
{{10'sd319, 11'sd839, 5'sd-10}, {13'sd2296, 13'sd2666, 11'sd921}, {12'sd-2010, 13'sd2684, 12'sd-1655}},
{{13'sd2599, 12'sd1869, 10'sd373}, {12'sd-1072, 12'sd1052, 12'sd-2047}, {12'sd1506, 12'sd1237, 10'sd-377}},
{{12'sd-1292, 11'sd-742, 11'sd-1023}, {10'sd294, 12'sd-1474, 12'sd1648}, {13'sd2227, 12'sd-1577, 13'sd-2877}},
{{13'sd-2429, 11'sd618, 11'sd-795}, {12'sd1893, 11'sd-886, 12'sd1849}, {13'sd-2058, 11'sd-771, 11'sd638}},
{{11'sd1021, 12'sd1461, 13'sd2219}, {13'sd-3062, 10'sd-312, 12'sd1534}, {13'sd-2606, 11'sd677, 12'sd-1202}},
{{8'sd98, 12'sd-1633, 11'sd891}, {13'sd2360, 12'sd1599, 12'sd-1893}, {9'sd195, 13'sd2379, 12'sd1758}},
{{11'sd895, 11'sd-989, 13'sd-2603}, {10'sd-510, 9'sd128, 10'sd-425}, {12'sd-1980, 11'sd596, 9'sd-246}},
{{13'sd2207, 13'sd-2138, 10'sd-384}, {11'sd925, 12'sd1706, 11'sd-904}, {12'sd1641, 11'sd515, 13'sd-2049}},
{{10'sd314, 9'sd193, 13'sd-4026}, {12'sd-1355, 7'sd-63, 12'sd1809}, {14'sd4515, 14'sd4298, 12'sd2028}},
{{10'sd-345, 13'sd2755, 13'sd-2672}, {13'sd-2146, 12'sd-1144, 11'sd-616}, {12'sd1897, 12'sd1847, 8'sd-123}},
{{13'sd-3219, 9'sd183, 12'sd1279}, {13'sd-2464, 13'sd-2212, 10'sd402}, {12'sd-1868, 12'sd-1852, 12'sd1308}},
{{11'sd752, 9'sd187, 13'sd3199}, {12'sd1827, 12'sd1434, 13'sd-2472}, {12'sd1691, 13'sd-2115, 12'sd1878}},
{{10'sd-486, 12'sd1489, 13'sd-2048}, {13'sd-2124, 11'sd801, 12'sd-1344}, {13'sd-2804, 12'sd1998, 9'sd232}},
{{11'sd977, 11'sd1013, 12'sd1468}, {12'sd1705, 12'sd1262, 13'sd2529}, {12'sd-1635, 13'sd-2088, 12'sd-1389}},
{{13'sd-2763, 12'sd1365, 11'sd-904}, {9'sd-243, 12'sd1815, 12'sd1283}, {8'sd126, 12'sd1619, 13'sd2416}},
{{12'sd1902, 10'sd-493, 12'sd1407}, {12'sd-1434, 10'sd-483, 13'sd2681}, {12'sd-1468, 12'sd1177, 12'sd-1910}},
{{12'sd-1770, 11'sd-535, 12'sd1277}, {12'sd-1964, 11'sd-534, 9'sd-198}, {13'sd-2512, 11'sd-615, 13'sd3805}},
{{13'sd2383, 5'sd13, 12'sd1783}, {11'sd-890, 8'sd117, 11'sd-826}, {13'sd-2264, 12'sd1878, 12'sd1037}},
{{11'sd-619, 12'sd-1193, 7'sd63}, {11'sd806, 9'sd-157, 8'sd-109}, {11'sd-913, 13'sd3433, 13'sd3306}},
{{12'sd-1071, 13'sd-2187, 13'sd-2555}, {7'sd-60, 12'sd-1356, 11'sd843}, {12'sd1610, 11'sd734, 13'sd2391}},
{{12'sd1445, 12'sd1781, 7'sd-59}, {9'sd203, 13'sd-2284, 11'sd-993}, {12'sd-1109, 12'sd-1219, 8'sd-127}},
{{12'sd-1774, 12'sd-1165, 10'sd310}, {10'sd326, 7'sd41, 8'sd126}, {7'sd-56, 11'sd857, 9'sd219}},
{{10'sd-372, 12'sd1435, 11'sd776}, {12'sd1722, 11'sd803, 12'sd1565}, {12'sd1140, 13'sd-2214, 11'sd658}},
{{12'sd1821, 13'sd2888, 13'sd-2234}, {12'sd-1629, 13'sd-2697, 12'sd-1498}, {13'sd-2406, 11'sd-636, 11'sd586}},
{{12'sd1978, 12'sd1721, 13'sd2271}, {12'sd-1861, 13'sd2662, 12'sd-1197}, {11'sd-660, 12'sd1708, 6'sd-29}},
{{14'sd-7306, 13'sd-2827, 12'sd-1686}, {13'sd-3611, 12'sd-1343, 13'sd-3212}, {13'sd-3584, 14'sd-4478, 13'sd-3635}},
{{11'sd-816, 11'sd995, 12'sd-1574}, {12'sd-1714, 11'sd716, 11'sd-891}, {10'sd-481, 13'sd2671, 13'sd-2069}},
{{12'sd1846, 10'sd272, 11'sd964}, {12'sd-1777, 12'sd1069, 13'sd2690}, {10'sd265, 13'sd-2857, 12'sd-1404}},
{{12'sd1160, 11'sd978, 13'sd3308}, {11'sd-845, 12'sd-1159, 12'sd1095}, {13'sd2608, 7'sd-51, 11'sd-606}},
{{11'sd-518, 12'sd2033, 12'sd-1841}, {12'sd1792, 13'sd2288, 11'sd-846}, {13'sd2684, 12'sd1932, 11'sd975}},
{{10'sd-499, 13'sd-2339, 7'sd-36}, {13'sd2062, 13'sd-2818, 12'sd1736}, {13'sd3178, 12'sd1567, 9'sd-143}},
{{13'sd2291, 11'sd946, 14'sd4730}, {13'sd2858, 11'sd808, 13'sd2457}, {13'sd-2967, 10'sd-455, 12'sd1831}},
{{10'sd-434, 12'sd-1299, 11'sd-989}, {11'sd685, 13'sd2962, 12'sd1507}, {11'sd-666, 10'sd264, 11'sd712}},
{{12'sd1065, 13'sd-2059, 13'sd-2247}, {12'sd-1913, 13'sd2445, 11'sd-568}, {11'sd-571, 13'sd-2992, 10'sd279}},
{{12'sd1667, 11'sd771, 13'sd-2720}, {13'sd-3125, 11'sd-586, 12'sd1869}, {13'sd-3960, 11'sd1008, 13'sd-2619}},
{{10'sd-281, 10'sd-405, 9'sd-188}, {11'sd953, 12'sd1750, 12'sd2001}, {11'sd-733, 10'sd-487, 11'sd-1002}},
{{12'sd1876, 12'sd1689, 11'sd829}, {12'sd1981, 8'sd-126, 11'sd733}, {12'sd-1629, 12'sd1556, 13'sd-2940}},
{{12'sd-1520, 13'sd-2660, 12'sd1345}, {13'sd2902, 12'sd1506, 9'sd183}, {10'sd-377, 13'sd-2614, 12'sd1234}},
{{13'sd-2697, 10'sd263, 12'sd-1737}, {13'sd-3159, 13'sd-2845, 14'sd-4393}, {15'sd-8334, 13'sd-3772, 14'sd-4325}},
{{13'sd-2363, 13'sd2467, 12'sd1809}, {10'sd-333, 11'sd765, 13'sd2371}, {13'sd2120, 12'sd1561, 12'sd-1599}},
{{12'sd1526, 12'sd-1802, 13'sd2350}, {12'sd1107, 13'sd2611, 12'sd-1767}, {11'sd682, 11'sd797, 11'sd972}},
{{12'sd2031, 11'sd685, 11'sd843}, {13'sd3452, 13'sd2740, 12'sd-1394}, {13'sd4070, 10'sd292, 13'sd2726}},
{{11'sd996, 12'sd-1238, 12'sd-1413}, {13'sd-2049, 13'sd2105, 11'sd911}, {11'sd923, 12'sd-1981, 9'sd-247}},
{{11'sd-942, 12'sd-1224, 13'sd2071}, {12'sd-1493, 11'sd-592, 12'sd1293}, {11'sd-872, 10'sd448, 9'sd218}},
{{12'sd1695, 11'sd514, 11'sd-1014}, {11'sd-871, 13'sd-2581, 10'sd373}, {13'sd-2349, 11'sd1006, 13'sd2266}},
{{11'sd-558, 11'sd-1004, 12'sd-1263}, {12'sd1537, 12'sd1904, 13'sd-2759}, {11'sd-745, 12'sd2028, 13'sd-2360}}},
{
{{12'sd1247, 13'sd2294, 12'sd-1576}, {11'sd987, 12'sd1863, 8'sd108}, {12'sd1807, 12'sd1953, 12'sd1382}},
{{10'sd403, 12'sd-1865, 13'sd2168}, {12'sd1393, 5'sd-12, 12'sd-1674}, {13'sd2757, 12'sd-1116, 5'sd-14}},
{{13'sd-3349, 11'sd-990, 13'sd2512}, {13'sd-2114, 13'sd2075, 11'sd-758}, {11'sd870, 13'sd2148, 12'sd-1719}},
{{13'sd-2488, 12'sd1450, 11'sd-990}, {12'sd-1689, 12'sd1039, 9'sd-238}, {12'sd-1326, 8'sd-126, 13'sd-2446}},
{{10'sd-328, 12'sd-1103, 14'sd5652}, {12'sd1150, 14'sd5986, 14'sd6921}, {10'sd-352, 14'sd4304, 14'sd5339}},
{{13'sd2424, 13'sd2178, 12'sd1412}, {10'sd-277, 13'sd2650, 10'sd325}, {12'sd1029, 10'sd-354, 13'sd2211}},
{{13'sd2513, 11'sd849, 14'sd4160}, {12'sd1991, 13'sd-3790, 12'sd1835}, {14'sd-4537, 13'sd-3672, 13'sd-2775}},
{{11'sd640, 11'sd-562, 13'sd-2273}, {12'sd-2002, 11'sd-587, 13'sd-2202}, {11'sd-747, 11'sd600, 10'sd-331}},
{{12'sd1822, 10'sd425, 10'sd-479}, {12'sd1469, 12'sd1762, 10'sd396}, {11'sd971, 11'sd-792, 13'sd3379}},
{{11'sd892, 12'sd1198, 13'sd3003}, {11'sd536, 8'sd96, 13'sd2716}, {12'sd1120, 12'sd1346, 9'sd201}},
{{13'sd-3539, 11'sd956, 13'sd-3364}, {13'sd-2626, 7'sd39, 13'sd-2491}, {14'sd-4440, 12'sd1081, 13'sd-2968}},
{{12'sd1671, 12'sd1930, 13'sd2428}, {10'sd352, 13'sd2877, 12'sd-1722}, {12'sd2027, 10'sd-371, 13'sd3209}},
{{10'sd398, 13'sd2675, 8'sd-96}, {13'sd2776, 12'sd-1584, 12'sd1950}, {10'sd297, 13'sd-2224, 13'sd3354}},
{{11'sd763, 11'sd-587, 13'sd-2404}, {12'sd1152, 13'sd-3064, 12'sd-1148}, {10'sd330, 11'sd782, 12'sd-1280}},
{{9'sd-232, 12'sd1535, 14'sd4657}, {12'sd-1645, 10'sd267, 11'sd-867}, {12'sd1109, 12'sd-1968, 13'sd-3029}},
{{9'sd-247, 7'sd-53, 11'sd-917}, {10'sd-296, 13'sd2529, 12'sd-1387}, {13'sd2112, 13'sd2495, 11'sd874}},
{{12'sd1268, 12'sd-1542, 12'sd1702}, {12'sd-1554, 9'sd198, 12'sd-1982}, {13'sd2730, 10'sd260, 13'sd-2262}},
{{13'sd-2729, 12'sd-1572, 13'sd3300}, {13'sd2389, 7'sd-44, 13'sd3612}, {12'sd-1605, 12'sd-1323, 13'sd3717}},
{{13'sd2403, 7'sd32, 11'sd-592}, {9'sd-242, 12'sd1062, 12'sd1588}, {11'sd672, 9'sd-143, 12'sd-1088}},
{{13'sd2886, 13'sd2072, 9'sd-168}, {12'sd-1146, 12'sd-1537, 12'sd1070}, {10'sd-480, 11'sd822, 13'sd-3276}},
{{12'sd1161, 12'sd-1414, 13'sd-2590}, {12'sd-2022, 10'sd510, 13'sd-2770}, {12'sd-1048, 13'sd-2814, 12'sd-1920}},
{{11'sd1016, 13'sd2072, 12'sd2029}, {12'sd1154, 9'sd182, 10'sd-369}, {13'sd2116, 13'sd2810, 12'sd1537}},
{{9'sd245, 11'sd967, 12'sd-1553}, {10'sd-269, 11'sd515, 12'sd-1040}, {12'sd-1097, 12'sd1328, 12'sd1262}},
{{12'sd1276, 13'sd-2285, 12'sd-1759}, {12'sd1755, 11'sd-987, 12'sd1410}, {12'sd-1535, 12'sd1381, 13'sd-2743}},
{{10'sd505, 11'sd-666, 12'sd1490}, {12'sd2009, 8'sd-73, 13'sd-2234}, {12'sd1273, 11'sd-532, 13'sd-2554}},
{{12'sd-1032, 12'sd1843, 13'sd3035}, {7'sd-46, 12'sd2037, 10'sd-347}, {12'sd-1551, 13'sd-2308, 9'sd251}},
{{14'sd-7240, 14'sd-7031, 14'sd-6127}, {13'sd-2699, 14'sd-7053, 12'sd-1851}, {13'sd-2791, 14'sd-4553, 11'sd-875}},
{{9'sd161, 12'sd-1912, 7'sd-53}, {9'sd-130, 13'sd2486, 13'sd2840}, {10'sd-419, 12'sd1447, 11'sd-791}},
{{12'sd-2040, 13'sd-3706, 12'sd-1391}, {14'sd-4661, 8'sd123, 11'sd520}, {12'sd-1416, 13'sd-3309, 13'sd-2183}},
{{12'sd-2018, 12'sd-1313, 12'sd1250}, {12'sd-1860, 12'sd1141, 12'sd-1212}, {11'sd-823, 13'sd-3076, 6'sd-21}},
{{12'sd1770, 12'sd1358, 12'sd-1093}, {8'sd103, 12'sd1763, 13'sd-2636}, {10'sd-494, 13'sd2637, 11'sd598}},
{{12'sd2043, 12'sd1097, 13'sd-2292}, {12'sd1370, 13'sd2133, 12'sd-1660}, {9'sd204, 12'sd-1877, 10'sd-508}},
{{10'sd344, 11'sd-708, 12'sd1543}, {11'sd794, 12'sd1604, 12'sd1993}, {13'sd2975, 11'sd1003, 12'sd-1852}},
{{13'sd-2483, 9'sd224, 11'sd-586}, {13'sd2080, 13'sd-2626, 12'sd-1459}, {13'sd-2181, 11'sd-787, 9'sd237}},
{{12'sd1986, 12'sd-2044, 11'sd-658}, {11'sd800, 12'sd1461, 10'sd-386}, {13'sd2573, 8'sd70, 10'sd-315}},
{{11'sd-888, 13'sd-2482, 7'sd-53}, {5'sd-8, 10'sd-492, 10'sd-384}, {11'sd597, 13'sd-3069, 13'sd-2102}},
{{11'sd596, 12'sd-1818, 12'sd-1181}, {8'sd123, 7'sd-59, 13'sd-2571}, {12'sd1051, 11'sd726, 13'sd-2861}},
{{12'sd1968, 13'sd2614, 12'sd1650}, {13'sd2373, 11'sd575, 9'sd229}, {13'sd-2123, 9'sd-198, 8'sd-80}},
{{13'sd2465, 12'sd-1806, 8'sd99}, {12'sd-1944, 12'sd1660, 12'sd1595}, {11'sd545, 12'sd-1491, 12'sd-1467}},
{{13'sd2055, 13'sd2951, 13'sd3067}, {11'sd922, 13'sd2186, 11'sd-988}, {10'sd267, 11'sd980, 12'sd-1832}},
{{6'sd-22, 13'sd2393, 11'sd-765}, {12'sd1501, 13'sd2522, 13'sd3858}, {11'sd670, 12'sd-1832, 12'sd-1320}},
{{13'sd2998, 13'sd2394, 13'sd3449}, {4'sd-6, 12'sd1948, 13'sd3699}, {13'sd-2240, 11'sd-806, 11'sd-969}},
{{14'sd-5466, 12'sd-1576, 7'sd52}, {14'sd-6331, 13'sd-2131, 13'sd-2540}, {13'sd-3347, 14'sd-5180, 14'sd-5720}},
{{14'sd-4630, 13'sd-3430, 11'sd-989}, {12'sd-1096, 12'sd-1068, 12'sd1105}, {13'sd-2443, 9'sd-178, 14'sd4338}},
{{10'sd-404, 11'sd562, 13'sd-2258}, {12'sd-1313, 11'sd832, 13'sd2109}, {13'sd-2616, 12'sd-1895, 12'sd-1890}},
{{13'sd2526, 10'sd279, 12'sd1143}, {12'sd1484, 13'sd2736, 11'sd918}, {11'sd967, 10'sd297, 8'sd-110}},
{{11'sd859, 13'sd2295, 13'sd-3331}, {9'sd-153, 12'sd-1827, 13'sd-3639}, {9'sd192, 12'sd-1139, 13'sd-2376}},
{{9'sd-248, 11'sd983, 11'sd-905}, {10'sd-422, 13'sd-2417, 12'sd1205}, {12'sd1805, 10'sd376, 13'sd-2391}},
{{12'sd1391, 8'sd-85, 13'sd-3027}, {9'sd-220, 12'sd-1737, 13'sd-3402}, {11'sd745, 13'sd-2614, 13'sd-3484}},
{{14'sd5597, 14'sd4779, 8'sd-93}, {14'sd4438, 14'sd4534, 10'sd-383}, {13'sd2323, 13'sd2964, 12'sd-1194}},
{{11'sd783, 12'sd-1743, 12'sd1309}, {13'sd-2111, 11'sd-753, 10'sd273}, {13'sd2057, 12'sd-1954, 12'sd-1449}},
{{13'sd-2944, 12'sd-1735, 11'sd926}, {13'sd2214, 10'sd438, 13'sd2735}, {11'sd-534, 13'sd2386, 13'sd2685}},
{{11'sd-908, 10'sd364, 12'sd1786}, {10'sd312, 13'sd2878, 12'sd-1596}, {11'sd-991, 12'sd-1832, 13'sd-3693}},
{{11'sd-654, 13'sd-3672, 9'sd-189}, {12'sd-1628, 12'sd-1062, 13'sd-2097}, {13'sd-2208, 8'sd126, 12'sd1364}},
{{13'sd3085, 11'sd856, 13'sd3794}, {10'sd-364, 11'sd931, 11'sd674}, {10'sd507, 13'sd-3824, 9'sd-140}},
{{13'sd2694, 10'sd-371, 13'sd-2881}, {11'sd769, 11'sd-765, 13'sd-2794}, {12'sd1878, 10'sd-315, 9'sd-201}},
{{13'sd-2072, 12'sd1230, 14'sd4591}, {13'sd2070, 13'sd3485, 13'sd2418}, {13'sd-3236, 11'sd-924, 11'sd-841}},
{{10'sd-286, 12'sd1084, 7'sd60}, {13'sd2096, 11'sd-551, 11'sd776}, {14'sd4312, 6'sd21, 9'sd-144}},
{{13'sd-2696, 12'sd1955, 9'sd-207}, {13'sd2525, 13'sd2174, 10'sd510}, {10'sd-268, 11'sd618, 11'sd729}},
{{10'sd388, 13'sd-2451, 12'sd1620}, {13'sd2286, 13'sd-2367, 11'sd559}, {10'sd506, 11'sd864, 8'sd-76}},
{{13'sd3091, 12'sd1545, 12'sd-2022}, {13'sd3498, 12'sd-1737, 12'sd-1996}, {11'sd996, 11'sd-533, 11'sd976}},
{{12'sd1204, 10'sd-428, 13'sd3127}, {12'sd1739, 9'sd-217, 13'sd2601}, {13'sd2250, 12'sd-1552, 10'sd-331}},
{{13'sd3022, 12'sd-1827, 11'sd556}, {13'sd3158, 12'sd-1668, 11'sd-792}, {12'sd1938, 13'sd2576, 12'sd-1703}},
{{12'sd-1971, 11'sd861, 13'sd-2401}, {14'sd-5524, 14'sd-5525, 10'sd278}, {12'sd-2031, 14'sd-4179, 13'sd-3502}}},
{
{{11'sd-751, 10'sd-290, 11'sd-576}, {12'sd1543, 12'sd-1715, 12'sd-1157}, {12'sd-1684, 12'sd-1885, 12'sd1527}},
{{11'sd620, 6'sd-29, 11'sd996}, {8'sd-65, 12'sd-1582, 11'sd-668}, {11'sd-773, 11'sd-955, 12'sd-1567}},
{{13'sd-2685, 13'sd2261, 13'sd-2319}, {13'sd-2054, 13'sd2680, 12'sd-1377}, {8'sd76, 12'sd1439, 13'sd-2684}},
{{13'sd2711, 13'sd-2399, 13'sd2612}, {13'sd-2248, 10'sd468, 13'sd2291}, {12'sd1293, 13'sd-2867, 11'sd-953}},
{{10'sd437, 13'sd2073, 12'sd1027}, {10'sd345, 11'sd-564, 11'sd889}, {10'sd-389, 10'sd258, 11'sd-737}},
{{11'sd-764, 12'sd1825, 13'sd-3852}, {12'sd-1168, 12'sd1308, 12'sd-1845}, {11'sd-581, 12'sd-1051, 13'sd-2103}},
{{13'sd3263, 13'sd3100, 12'sd1445}, {13'sd3133, 12'sd1517, 13'sd-3981}, {7'sd61, 12'sd-1841, 10'sd-276}},
{{13'sd2783, 11'sd722, 12'sd1456}, {12'sd1928, 12'sd1852, 12'sd-1809}, {12'sd-1967, 9'sd-193, 11'sd940}},
{{12'sd-1258, 12'sd1886, 11'sd-860}, {12'sd-1438, 8'sd-74, 12'sd1545}, {13'sd2295, 12'sd-1441, 6'sd-19}},
{{13'sd2187, 12'sd-1490, 12'sd1669}, {13'sd2292, 10'sd403, 12'sd-1473}, {5'sd12, 13'sd-2653, 11'sd-859}},
{{12'sd-1140, 13'sd-2268, 12'sd-1883}, {12'sd-2032, 11'sd-1011, 13'sd-2606}, {12'sd-1481, 12'sd-1511, 11'sd-993}},
{{8'sd-66, 13'sd2349, 7'sd-61}, {12'sd2011, 13'sd-2197, 12'sd1196}, {13'sd2341, 12'sd1608, 12'sd1501}},
{{13'sd2290, 13'sd3088, 12'sd-1253}, {12'sd-1390, 13'sd2639, 12'sd-1474}, {10'sd-267, 12'sd1630, 12'sd-1287}},
{{11'sd-956, 13'sd2572, 10'sd-366}, {12'sd-1416, 12'sd-1609, 12'sd1623}, {12'sd1503, 11'sd903, 13'sd-2081}},
{{13'sd-3220, 11'sd-874, 13'sd-2503}, {12'sd-1720, 12'sd1100, 13'sd-2652}, {12'sd-1223, 13'sd4058, 11'sd-778}},
{{12'sd1614, 12'sd1929, 12'sd-1248}, {12'sd-1653, 13'sd2337, 13'sd2158}, {13'sd-2438, 13'sd2886, 12'sd-1034}},
{{13'sd-2138, 13'sd-2727, 12'sd1468}, {12'sd-1420, 12'sd-1332, 12'sd-1967}, {10'sd-465, 13'sd-2518, 10'sd-295}},
{{12'sd1573, 13'sd-2286, 12'sd1321}, {10'sd-423, 13'sd-2488, 11'sd-641}, {12'sd1960, 12'sd1886, 12'sd-1833}},
{{12'sd1026, 12'sd-1840, 13'sd2056}, {13'sd-2564, 12'sd-1223, 10'sd-498}, {12'sd-1184, 11'sd-599, 10'sd339}},
{{11'sd932, 9'sd-153, 12'sd1778}, {12'sd1994, 13'sd-2402, 12'sd-1308}, {9'sd-246, 12'sd-1821, 12'sd1279}},
{{12'sd-1212, 12'sd2001, 13'sd-2339}, {12'sd1318, 11'sd-761, 13'sd2449}, {12'sd1304, 10'sd409, 12'sd1278}},
{{11'sd724, 12'sd1967, 13'sd2645}, {13'sd-2525, 12'sd1866, 10'sd380}, {12'sd1338, 12'sd1058, 13'sd2154}},
{{10'sd497, 10'sd-407, 13'sd2048}, {11'sd-790, 10'sd-260, 13'sd2729}, {12'sd-1334, 12'sd-1723, 12'sd1721}},
{{9'sd-157, 12'sd-1383, 13'sd-2216}, {11'sd-661, 12'sd-1309, 13'sd-2384}, {13'sd-2582, 12'sd1610, 10'sd423}},
{{13'sd2187, 12'sd-1542, 12'sd-1067}, {13'sd2106, 11'sd897, 12'sd1170}, {12'sd-1368, 11'sd-700, 11'sd695}},
{{13'sd-2384, 10'sd256, 12'sd1805}, {13'sd2397, 10'sd423, 12'sd-2032}, {12'sd-1370, 11'sd544, 13'sd2575}},
{{13'sd3592, 13'sd-2837, 13'sd-3937}, {12'sd1522, 12'sd-2037, 14'sd-4205}, {13'sd2602, 10'sd-319, 12'sd-1593}},
{{8'sd66, 11'sd989, 10'sd459}, {12'sd-1086, 10'sd311, 10'sd314}, {9'sd-158, 10'sd-351, 12'sd-2035}},
{{12'sd-1256, 13'sd2448, 12'sd-1303}, {10'sd-271, 13'sd-2243, 13'sd-2162}, {11'sd942, 12'sd1287, 13'sd-2363}},
{{8'sd118, 11'sd926, 11'sd884}, {13'sd-2913, 11'sd728, 13'sd-2275}, {12'sd-1544, 12'sd1811, 10'sd320}},
{{12'sd-1775, 13'sd-2105, 9'sd252}, {11'sd-656, 13'sd2238, 9'sd132}, {13'sd2567, 10'sd-404, 12'sd-1525}},
{{10'sd-290, 13'sd-2174, 12'sd-1784}, {12'sd-1397, 10'sd317, 12'sd-1742}, {12'sd1217, 10'sd306, 11'sd-895}},
{{13'sd3044, 12'sd1755, 11'sd940}, {9'sd-255, 12'sd-1713, 13'sd-2122}, {13'sd2586, 11'sd915, 13'sd2195}},
{{12'sd1475, 12'sd-1596, 10'sd335}, {12'sd-1436, 12'sd1266, 13'sd-2073}, {12'sd1170, 12'sd-1653, 12'sd1891}},
{{12'sd1198, 12'sd-1844, 12'sd1374}, {10'sd337, 12'sd-1812, 13'sd2596}, {12'sd1540, 13'sd2365, 12'sd1118}},
{{11'sd673, 12'sd1772, 12'sd1483}, {12'sd1277, 12'sd-1032, 12'sd-1158}, {13'sd-2070, 13'sd2768, 12'sd1185}},
{{13'sd2900, 13'sd-2165, 11'sd-726}, {13'sd2542, 13'sd3091, 13'sd3244}, {11'sd647, 12'sd-1125, 12'sd1651}},
{{9'sd137, 12'sd-1396, 13'sd2484}, {13'sd3148, 12'sd1839, 12'sd1307}, {10'sd-365, 13'sd-2288, 10'sd-488}},
{{11'sd967, 12'sd1880, 13'sd-2868}, {12'sd-1981, 12'sd-1153, 11'sd-777}, {13'sd-2616, 12'sd1256, 12'sd-1829}},
{{12'sd1463, 11'sd-866, 11'sd-906}, {13'sd-2542, 11'sd1006, 10'sd-462}, {10'sd-443, 12'sd1294, 12'sd-1150}},
{{13'sd2164, 11'sd981, 12'sd-1989}, {11'sd-844, 12'sd1716, 11'sd-978}, {13'sd2668, 12'sd1229, 12'sd-1439}},
{{9'sd195, 11'sd846, 11'sd796}, {13'sd2368, 12'sd1536, 13'sd2164}, {12'sd1735, 12'sd1439, 12'sd1112}},
{{13'sd-3786, 11'sd-757, 12'sd1994}, {12'sd1166, 12'sd1458, 12'sd1309}, {12'sd-1840, 7'sd-43, 13'sd-2283}},
{{11'sd-932, 14'sd-4754, 13'sd-3957}, {9'sd-172, 9'sd-144, 13'sd-2234}, {14'sd6999, 14'sd4224, 12'sd-1795}},
{{10'sd-338, 12'sd2005, 12'sd-1772}, {13'sd2536, 12'sd1211, 11'sd-765}, {12'sd-1446, 11'sd944, 13'sd-2056}},
{{12'sd1208, 12'sd1712, 13'sd-2398}, {12'sd2025, 12'sd1098, 12'sd-1743}, {12'sd1817, 10'sd430, 12'sd1130}},
{{12'sd-1722, 12'sd-1071, 10'sd-264}, {12'sd-1192, 13'sd-2442, 13'sd-2102}, {11'sd899, 12'sd-1637, 11'sd-766}},
{{11'sd-992, 11'sd910, 12'sd-1710}, {12'sd-1979, 12'sd-1791, 13'sd-2240}, {12'sd1744, 13'sd2468, 13'sd3185}},
{{11'sd934, 10'sd-438, 12'sd1192}, {11'sd-714, 11'sd932, 12'sd-1426}, {13'sd-2221, 13'sd-2212, 11'sd-758}},
{{13'sd2900, 12'sd-1608, 14'sd4248}, {11'sd691, 12'sd1215, 13'sd2365}, {12'sd-1355, 12'sd-1225, 12'sd1921}},
{{10'sd483, 10'sd-491, 13'sd2283}, {12'sd-1056, 10'sd447, 10'sd485}, {12'sd1714, 12'sd1888, 12'sd-1590}},
{{13'sd-2093, 12'sd2006, 12'sd-2031}, {12'sd1548, 13'sd2087, 11'sd-682}, {12'sd-1885, 11'sd629, 12'sd-1200}},
{{10'sd-448, 10'sd412, 13'sd-2308}, {13'sd-2439, 11'sd555, 11'sd-698}, {8'sd-101, 13'sd2508, 11'sd610}},
{{12'sd1515, 11'sd-861, 10'sd356}, {13'sd2466, 8'sd76, 12'sd-1475}, {11'sd550, 13'sd-2090, 12'sd1746}},
{{10'sd-443, 11'sd819, 12'sd-1657}, {10'sd-432, 11'sd658, 11'sd622}, {10'sd-267, 13'sd-3480, 12'sd-1670}},
{{12'sd-1888, 13'sd-2947, 8'sd106}, {13'sd2171, 7'sd45, 10'sd-264}, {10'sd-446, 13'sd-2127, 12'sd1233}},
{{14'sd4334, 12'sd1629, 14'sd5037}, {13'sd2887, 10'sd260, 13'sd3491}, {13'sd-3277, 11'sd942, 12'sd-1371}},
{{9'sd157, 12'sd1643, 11'sd536}, {8'sd-123, 9'sd164, 13'sd2125}, {10'sd-492, 13'sd2306, 12'sd1641}},
{{12'sd1051, 12'sd1370, 12'sd1640}, {11'sd580, 9'sd254, 12'sd-1276}, {12'sd1520, 9'sd189, 13'sd2048}},
{{11'sd-583, 13'sd2208, 12'sd-1330}, {12'sd-1094, 13'sd2364, 12'sd-1796}, {13'sd-3187, 11'sd885, 13'sd-2386}},
{{11'sd-542, 12'sd1638, 13'sd-2073}, {10'sd-274, 12'sd-1210, 12'sd1725}, {13'sd2382, 12'sd-1444, 12'sd1779}},
{{10'sd491, 7'sd52, 9'sd-211}, {12'sd-1526, 12'sd1387, 11'sd-856}, {13'sd-3055, 10'sd459, 10'sd-350}},
{{13'sd4053, 12'sd-2027, 12'sd-1524}, {13'sd2954, 11'sd-617, 13'sd2409}, {12'sd-1898, 8'sd88, 12'sd1909}},
{{13'sd-3482, 13'sd-3131, 12'sd-1493}, {11'sd577, 5'sd12, 13'sd-2521}, {13'sd-2431, 12'sd-1919, 10'sd285}}},
{
{{13'sd-2051, 12'sd-1297, 11'sd-869}, {13'sd-2072, 11'sd1009, 13'sd2398}, {12'sd-1712, 13'sd-2525, 9'sd-138}},
{{12'sd-1158, 12'sd-1493, 12'sd1383}, {12'sd-1905, 13'sd-2886, 13'sd-2697}, {12'sd-1878, 13'sd-3321, 11'sd912}},
{{12'sd1089, 10'sd423, 8'sd-66}, {11'sd-530, 12'sd1139, 13'sd-2083}, {9'sd203, 12'sd1282, 9'sd132}},
{{13'sd2699, 12'sd1780, 12'sd1194}, {11'sd660, 10'sd-292, 12'sd-1663}, {12'sd1301, 12'sd-1325, 8'sd96}},
{{13'sd-2066, 12'sd-1106, 13'sd-3999}, {11'sd-963, 10'sd-432, 12'sd-1873}, {12'sd-1076, 12'sd-1314, 9'sd-146}},
{{10'sd-433, 13'sd-2157, 13'sd-2195}, {13'sd-2197, 13'sd-2132, 12'sd-1281}, {12'sd-2031, 10'sd364, 13'sd-2723}},
{{12'sd-1245, 13'sd-2431, 12'sd1206}, {13'sd3059, 11'sd536, 11'sd-537}, {14'sd4463, 10'sd502, 12'sd1954}},
{{12'sd-1444, 13'sd-2652, 10'sd287}, {13'sd-2268, 11'sd562, 11'sd-867}, {9'sd211, 11'sd-708, 11'sd737}},
{{12'sd-1378, 10'sd-462, 13'sd2506}, {11'sd-523, 11'sd862, 11'sd984}, {5'sd-10, 11'sd-912, 12'sd1157}},
{{13'sd2149, 11'sd838, 12'sd-1651}, {12'sd-1775, 11'sd1020, 11'sd-984}, {12'sd-1114, 13'sd2573, 13'sd-2191}},
{{11'sd529, 13'sd2412, 11'sd-960}, {13'sd2767, 12'sd1487, 11'sd-542}, {12'sd2022, 9'sd-192, 13'sd2445}},
{{12'sd-1301, 9'sd-199, 12'sd-1747}, {12'sd-1120, 13'sd-3033, 10'sd-399}, {12'sd1935, 9'sd-175, 12'sd-1386}},
{{13'sd-2284, 13'sd-2747, 13'sd-2258}, {12'sd-1721, 11'sd870, 12'sd1803}, {13'sd-2294, 11'sd-920, 12'sd-1683}},
{{13'sd2598, 13'sd2496, 12'sd-1954}, {12'sd1356, 11'sd-734, 11'sd681}, {13'sd-2895, 12'sd1332, 12'sd1969}},
{{9'sd-174, 13'sd3285, 13'sd3656}, {13'sd2175, 11'sd528, 13'sd2956}, {12'sd1424, 12'sd-1194, 12'sd-1496}},
{{12'sd1597, 12'sd1501, 10'sd462}, {10'sd-434, 13'sd-2454, 12'sd-1150}, {12'sd-1533, 11'sd-668, 10'sd327}},
{{11'sd670, 13'sd2210, 13'sd2515}, {12'sd2034, 12'sd-2005, 11'sd-686}, {13'sd2349, 8'sd-95, 11'sd-556}},
{{13'sd-2185, 13'sd-2654, 13'sd-2907}, {13'sd-2373, 13'sd-2449, 12'sd-1287}, {12'sd1428, 13'sd2077, 7'sd46}},
{{13'sd2372, 13'sd2313, 10'sd-373}, {13'sd2775, 12'sd1780, 12'sd1865}, {12'sd-1076, 13'sd-2126, 12'sd-1123}},
{{12'sd-1561, 11'sd832, 12'sd1547}, {12'sd1148, 8'sd93, 5'sd-12}, {13'sd2475, 8'sd-89, 12'sd-1598}},
{{13'sd-2665, 12'sd1543, 13'sd-2545}, {11'sd-648, 13'sd2692, 12'sd-1298}, {12'sd1784, 12'sd1454, 10'sd-392}},
{{13'sd-2697, 12'sd1369, 12'sd1953}, {13'sd-2562, 10'sd349, 12'sd1667}, {10'sd439, 11'sd-858, 12'sd1744}},
{{13'sd-2864, 13'sd2081, 12'sd1364}, {13'sd-2073, 12'sd-1819, 11'sd-616}, {13'sd-2424, 11'sd-547, 6'sd-19}},
{{12'sd-1964, 13'sd2184, 12'sd-1323}, {10'sd-306, 9'sd-254, 4'sd-5}, {11'sd-977, 12'sd-1181, 10'sd346}},
{{13'sd2763, 13'sd2471, 11'sd-572}, {12'sd1797, 8'sd83, 13'sd2266}, {10'sd-449, 12'sd1189, 10'sd-440}},
{{13'sd2459, 13'sd-2490, 12'sd1432}, {13'sd2132, 13'sd2253, 13'sd-2645}, {13'sd-2121, 8'sd90, 12'sd-1258}},
{{13'sd2475, 11'sd889, 10'sd363}, {8'sd-66, 11'sd918, 9'sd130}, {13'sd3634, 13'sd2412, 9'sd-196}},
{{12'sd1870, 13'sd-2354, 12'sd1643}, {11'sd-673, 13'sd-2371, 11'sd854}, {12'sd1336, 13'sd3030, 9'sd236}},
{{13'sd2228, 11'sd-743, 9'sd-194}, {12'sd-1032, 12'sd-1674, 11'sd-1011}, {13'sd2574, 13'sd3053, 13'sd2500}},
{{12'sd-1263, 11'sd948, 11'sd-786}, {13'sd2896, 12'sd1885, 13'sd2391}, {12'sd1580, 13'sd3206, 12'sd1487}},
{{12'sd-1363, 10'sd-423, 11'sd-919}, {13'sd-2836, 13'sd-2299, 12'sd1770}, {12'sd-1804, 13'sd2442, 9'sd235}},
{{12'sd-1778, 12'sd-1398, 10'sd348}, {13'sd-2371, 12'sd-1577, 12'sd-1309}, {12'sd1927, 13'sd2311, 11'sd584}},
{{12'sd1621, 10'sd-305, 13'sd2196}, {12'sd-1553, 12'sd-1244, 13'sd-2505}, {11'sd710, 12'sd1849, 12'sd1381}},
{{12'sd1500, 13'sd2188, 13'sd3065}, {13'sd2577, 10'sd-338, 9'sd-175}, {12'sd1910, 11'sd-683, 13'sd3316}},
{{12'sd-2003, 11'sd-680, 10'sd300}, {13'sd-2867, 11'sd724, 13'sd2825}, {9'sd-191, 12'sd1094, 13'sd2706}},
{{13'sd2346, 13'sd-2146, 11'sd624}, {13'sd2907, 9'sd-184, 12'sd1095}, {13'sd2832, 13'sd-2205, 11'sd651}},
{{12'sd-1748, 11'sd-596, 12'sd1635}, {12'sd-1411, 13'sd3917, 13'sd2094}, {12'sd2046, 13'sd3287, 14'sd4461}},
{{11'sd-792, 10'sd-433, 12'sd-1121}, {12'sd-1601, 11'sd823, 9'sd133}, {12'sd1192, 13'sd2433, 11'sd-965}},
{{13'sd-2122, 9'sd200, 12'sd-1188}, {13'sd-2423, 11'sd-621, 13'sd2437}, {12'sd-1308, 13'sd2638, 13'sd2105}},
{{13'sd2420, 12'sd1555, 9'sd169}, {11'sd-584, 8'sd-91, 11'sd607}, {12'sd1132, 10'sd-306, 12'sd1564}},
{{12'sd2013, 13'sd-2808, 13'sd-2106}, {13'sd2084, 13'sd-2195, 11'sd-523}, {12'sd1572, 13'sd-2567, 12'sd-1787}},
{{9'sd-166, 10'sd-299, 10'sd-305}, {13'sd-2819, 13'sd-2381, 13'sd2291}, {12'sd-1510, 12'sd-1796, 9'sd-149}},
{{10'sd-271, 9'sd171, 13'sd-2216}, {12'sd1888, 12'sd1818, 13'sd3307}, {14'sd4901, 12'sd1358, 7'sd-43}},
{{12'sd1095, 13'sd-3190, 10'sd362}, {10'sd-294, 13'sd-2219, 11'sd-552}, {13'sd-3046, 13'sd-2292, 12'sd-1496}},
{{12'sd1971, 12'sd1359, 9'sd-212}, {13'sd2084, 8'sd102, 12'sd1533}, {13'sd-2478, 13'sd2533, 9'sd229}},
{{12'sd-1993, 10'sd-394, 12'sd-1073}, {12'sd-1161, 12'sd-1136, 13'sd2519}, {13'sd-2828, 12'sd-1290, 12'sd-1560}},
{{12'sd1662, 9'sd-207, 13'sd3006}, {13'sd-2556, 11'sd-759, 13'sd3582}, {10'sd477, 11'sd-921, 11'sd928}},
{{10'sd-289, 10'sd-331, 13'sd2458}, {12'sd1457, 12'sd1073, 13'sd2182}, {12'sd-1746, 9'sd-132, 11'sd994}},
{{13'sd2180, 12'sd-1292, 12'sd1175}, {12'sd-1441, 6'sd-27, 12'sd-1186}, {11'sd-843, 12'sd-1864, 13'sd2375}},
{{11'sd835, 12'sd1862, 12'sd1770}, {13'sd-3169, 10'sd357, 11'sd970}, {11'sd703, 13'sd2323, 13'sd2089}},
{{12'sd-1187, 10'sd433, 12'sd-1654}, {13'sd-2063, 11'sd-815, 10'sd-331}, {9'sd-220, 12'sd-1576, 10'sd269}},
{{12'sd1571, 12'sd-1618, 12'sd1837}, {13'sd-2440, 12'sd-1026, 12'sd1898}, {13'sd-2566, 12'sd1734, 8'sd-89}},
{{13'sd-2426, 12'sd-1951, 13'sd-2894}, {12'sd1570, 12'sd1858, 7'sd-32}, {13'sd3627, 13'sd3079, 13'sd2611}},
{{11'sd-1020, 12'sd1454, 11'sd-781}, {12'sd-1716, 12'sd1249, 7'sd61}, {12'sd-1885, 13'sd-2546, 10'sd475}},
{{13'sd-2167, 10'sd443, 12'sd1148}, {7'sd-60, 12'sd1388, 13'sd-3632}, {13'sd3974, 12'sd1213, 12'sd-2046}},
{{13'sd2650, 12'sd1173, 10'sd506}, {13'sd2817, 13'sd2809, 12'sd1413}, {12'sd-1306, 12'sd1889, 12'sd-1384}},
{{7'sd-60, 11'sd-753, 12'sd-1058}, {12'sd1731, 11'sd-752, 14'sd-4835}, {11'sd612, 12'sd1683, 12'sd1125}},
{{12'sd1031, 13'sd2122, 10'sd432}, {12'sd-1394, 12'sd-1963, 10'sd295}, {5'sd9, 12'sd1241, 12'sd-1330}},
{{11'sd-864, 12'sd-1885, 11'sd-935}, {12'sd1721, 11'sd986, 12'sd2039}, {9'sd-211, 12'sd-2038, 13'sd-2201}},
{{12'sd-1096, 12'sd1475, 12'sd1641}, {12'sd-1252, 13'sd2505, 12'sd-1925}, {11'sd730, 12'sd1102, 8'sd115}},
{{11'sd-742, 13'sd-2227, 10'sd316}, {12'sd-1466, 7'sd42, 11'sd727}, {13'sd-3229, 9'sd-242, 12'sd-1680}},
{{13'sd2077, 13'sd2349, 10'sd313}, {8'sd-100, 13'sd-2651, 12'sd-1270}, {12'sd-1694, 9'sd-216, 11'sd-886}},
{{12'sd1951, 12'sd-1473, 12'sd-1323}, {12'sd-1438, 13'sd2885, 12'sd1474}, {12'sd-1496, 9'sd-158, 13'sd-2852}},
{{12'sd-1413, 10'sd356, 12'sd1067}, {13'sd2884, 11'sd-830, 13'sd2172}, {13'sd2982, 9'sd-189, 4'sd-5}}},
{
{{12'sd-1233, 13'sd-2331, 12'sd-1660}, {13'sd-2806, 13'sd-3042, 13'sd2244}, {11'sd878, 8'sd-106, 12'sd1381}},
{{9'sd146, 13'sd2064, 12'sd-1767}, {10'sd-440, 11'sd-987, 12'sd-1529}, {11'sd743, 11'sd925, 9'sd-210}},
{{13'sd-2581, 11'sd861, 12'sd-1233}, {11'sd-816, 13'sd-2399, 7'sd-34}, {12'sd-1385, 12'sd1623, 13'sd-2521}},
{{12'sd-1580, 12'sd1984, 13'sd-2985}, {8'sd-97, 11'sd998, 12'sd-1959}, {12'sd-1131, 13'sd3249, 13'sd2713}},
{{13'sd2520, 13'sd2234, 11'sd-999}, {11'sd-622, 13'sd2493, 13'sd2488}, {8'sd67, 11'sd-949, 11'sd744}},
{{14'sd4119, 13'sd2468, 13'sd-2575}, {11'sd525, 12'sd1245, 14'sd-5126}, {11'sd-698, 8'sd74, 14'sd-4755}},
{{13'sd4040, 13'sd3426, 9'sd194}, {13'sd3244, 13'sd3572, 10'sd-316}, {13'sd3580, 13'sd3544, 13'sd2160}},
{{13'sd-2088, 11'sd-635, 13'sd2090}, {12'sd1313, 13'sd2051, 13'sd2147}, {13'sd2882, 11'sd756, 10'sd351}},
{{10'sd327, 13'sd2097, 9'sd216}, {12'sd-1254, 11'sd-633, 12'sd1713}, {12'sd1841, 12'sd-1543, 13'sd2143}},
{{12'sd-1732, 9'sd-182, 13'sd3193}, {12'sd1833, 12'sd1151, 13'sd2818}, {11'sd-1002, 12'sd1105, 11'sd-858}},
{{12'sd-1954, 12'sd1865, 10'sd-317}, {12'sd-1598, 10'sd-277, 12'sd-1124}, {13'sd-2856, 12'sd1637, 10'sd407}},
{{13'sd-2186, 12'sd1051, 12'sd1921}, {12'sd-1364, 12'sd1669, 13'sd-3444}, {12'sd1516, 11'sd-768, 12'sd-1699}},
{{11'sd-626, 12'sd1953, 13'sd2060}, {13'sd-2988, 12'sd-1397, 13'sd-2262}, {13'sd-2519, 12'sd1337, 10'sd-386}},
{{12'sd1217, 12'sd-1901, 8'sd79}, {13'sd-2423, 13'sd-2367, 13'sd2740}, {12'sd1402, 13'sd-2678, 13'sd3156}},
{{12'sd-1601, 13'sd-2426, 14'sd-4442}, {13'sd3851, 12'sd1503, 13'sd-2407}, {13'sd2471, 12'sd1765, 12'sd2001}},
{{12'sd-1043, 13'sd-2083, 13'sd-2320}, {9'sd205, 12'sd1445, 13'sd-2650}, {12'sd-1357, 13'sd-2442, 12'sd-1494}},
{{12'sd-1539, 12'sd-1898, 13'sd-2509}, {11'sd-575, 12'sd-1228, 12'sd1138}, {12'sd1490, 9'sd-222, 13'sd-2781}},
{{11'sd728, 10'sd-444, 12'sd-1395}, {12'sd1774, 12'sd1065, 13'sd2805}, {13'sd-2176, 13'sd2738, 12'sd-1052}},
{{12'sd2007, 13'sd-2287, 13'sd2890}, {13'sd2539, 12'sd-1942, 12'sd-2041}, {11'sd691, 13'sd-2143, 13'sd2881}},
{{12'sd-1893, 13'sd2998, 13'sd2461}, {13'sd-2215, 11'sd1012, 12'sd-1194}, {13'sd2500, 7'sd39, 13'sd2074}},
{{12'sd1350, 13'sd-2561, 10'sd362}, {8'sd-89, 12'sd1403, 10'sd362}, {10'sd274, 11'sd723, 10'sd500}},
{{11'sd824, 11'sd857, 13'sd-2400}, {12'sd1625, 11'sd-1010, 11'sd-711}, {12'sd-1565, 12'sd-1348, 12'sd1100}},
{{11'sd888, 11'sd-603, 13'sd-2512}, {12'sd-1700, 12'sd-2005, 12'sd-1710}, {12'sd1255, 13'sd-2095, 13'sd-2961}},
{{12'sd-1058, 12'sd-1485, 11'sd757}, {12'sd1394, 13'sd2483, 13'sd2385}, {12'sd-1118, 13'sd-2051, 11'sd-650}},
{{13'sd-2648, 12'sd1400, 13'sd-2325}, {13'sd-2428, 11'sd-882, 9'sd178}, {8'sd64, 10'sd259, 12'sd1380}},
{{13'sd-2135, 11'sd794, 13'sd-2084}, {13'sd-2423, 11'sd-694, 12'sd1386}, {10'sd-369, 12'sd1311, 13'sd-2359}},
{{12'sd-1443, 13'sd3527, 12'sd1872}, {13'sd-2392, 13'sd2674, 12'sd1217}, {11'sd-784, 13'sd2769, 13'sd2563}},
{{13'sd2433, 13'sd-2749, 12'sd-1360}, {12'sd-1245, 11'sd-823, 13'sd-2186}, {10'sd-490, 10'sd380, 12'sd-1029}},
{{13'sd-3549, 13'sd-2867, 13'sd-2621}, {13'sd-3027, 13'sd-3103, 12'sd1108}, {7'sd52, 11'sd-565, 12'sd-1155}},
{{10'sd485, 10'sd-317, 12'sd1900}, {13'sd2688, 11'sd-1004, 12'sd-1981}, {10'sd350, 12'sd1120, 9'sd-153}},
{{13'sd2382, 12'sd-1587, 10'sd-477}, {13'sd2273, 13'sd-2735, 12'sd-1435}, {13'sd-2260, 8'sd97, 11'sd-899}},
{{10'sd350, 9'sd205, 11'sd1016}, {13'sd-2209, 12'sd1577, 10'sd-487}, {7'sd-59, 13'sd-2278, 13'sd-2449}},
{{8'sd105, 12'sd1459, 11'sd-542}, {12'sd1254, 10'sd-488, 10'sd371}, {13'sd-2394, 12'sd-1547, 6'sd22}},
{{12'sd1209, 12'sd1158, 11'sd644}, {11'sd845, 13'sd-2483, 12'sd-1919}, {12'sd1814, 9'sd-133, 9'sd168}},
{{12'sd1378, 9'sd170, 12'sd2045}, {13'sd4047, 13'sd-2673, 10'sd358}, {11'sd596, 11'sd-936, 13'sd-3179}},
{{13'sd-2162, 12'sd-1053, 13'sd-3173}, {10'sd-294, 11'sd646, 12'sd-1901}, {13'sd-2217, 10'sd-286, 12'sd-1897}},
{{13'sd-2078, 13'sd-2661, 5'sd-10}, {13'sd3353, 12'sd2031, 12'sd1459}, {12'sd1409, 6'sd-19, 13'sd-4090}},
{{12'sd1292, 8'sd100, 12'sd-2029}, {12'sd1663, 13'sd3127, 10'sd485}, {12'sd1502, 11'sd1000, 11'sd659}},
{{11'sd744, 8'sd117, 7'sd-32}, {12'sd1610, 10'sd444, 10'sd408}, {11'sd-801, 12'sd-1314, 12'sd-1072}},
{{13'sd-2225, 13'sd2344, 13'sd-2814}, {11'sd-911, 13'sd-2580, 13'sd-2495}, {11'sd-971, 12'sd1603, 13'sd-2602}},
{{7'sd38, 13'sd3451, 9'sd-212}, {12'sd1294, 11'sd-832, 10'sd-352}, {9'sd-159, 13'sd2607, 11'sd611}},
{{13'sd-2310, 13'sd-3300, 8'sd-93}, {11'sd928, 11'sd994, 12'sd1820}, {12'sd1942, 11'sd-883, 12'sd1533}},
{{11'sd837, 13'sd-3572, 12'sd-1549}, {11'sd543, 12'sd-1527, 13'sd2434}, {10'sd-341, 11'sd-734, 11'sd-993}},
{{14'sd-7451, 14'sd-5729, 12'sd-1967}, {13'sd-2586, 12'sd1688, 13'sd-3317}, {13'sd-3165, 13'sd-2462, 13'sd-3759}},
{{11'sd935, 13'sd2847, 12'sd-1913}, {11'sd645, 13'sd-2182, 11'sd-873}, {11'sd802, 12'sd1762, 11'sd831}},
{{12'sd1764, 13'sd-3249, 13'sd-2433}, {11'sd882, 12'sd1233, 13'sd-3758}, {11'sd1021, 11'sd-642, 13'sd-3723}},
{{12'sd-1105, 12'sd1968, 13'sd2453}, {12'sd-1181, 10'sd-269, 13'sd-2417}, {12'sd1748, 13'sd2150, 11'sd787}},
{{12'sd1212, 13'sd-2334, 12'sd-1597}, {10'sd510, 12'sd1306, 13'sd2817}, {13'sd2721, 13'sd-2320, 12'sd-1176}},
{{12'sd-1258, 11'sd941, 13'sd-2916}, {11'sd-637, 13'sd-2231, 10'sd-407}, {14'sd4780, 13'sd2179, 11'sd780}},
{{14'sd4435, 6'sd31, 12'sd1558}, {12'sd1762, 12'sd-1600, 12'sd1219}, {10'sd-287, 9'sd134, 12'sd1440}},
{{13'sd3673, 12'sd1840, 13'sd3314}, {13'sd2509, 13'sd-2508, 8'sd90}, {13'sd-2133, 11'sd-588, 9'sd-205}},
{{12'sd-1540, 13'sd2561, 11'sd-1003}, {13'sd-2142, 11'sd707, 13'sd2085}, {11'sd745, 11'sd585, 11'sd620}},
{{13'sd-3936, 11'sd-927, 12'sd1189}, {11'sd-869, 12'sd1498, 11'sd-536}, {12'sd1175, 11'sd817, 5'sd-13}},
{{13'sd-2273, 12'sd1534, 12'sd2002}, {12'sd-2019, 12'sd-1518, 12'sd-1415}, {12'sd-1983, 11'sd-594, 11'sd-915}},
{{12'sd-1299, 12'sd-1094, 10'sd-392}, {13'sd3628, 12'sd1834, 12'sd-1682}, {13'sd3556, 13'sd2124, 13'sd2843}},
{{12'sd1961, 11'sd687, 13'sd-3244}, {11'sd-945, 10'sd-333, 12'sd-1735}, {12'sd-1783, 12'sd1794, 12'sd1161}},
{{7'sd46, 11'sd547, 12'sd1710}, {11'sd896, 14'sd4389, 14'sd4626}, {7'sd-39, 11'sd961, 14'sd4799}},
{{13'sd2051, 12'sd1468, 12'sd2033}, {12'sd-1566, 12'sd-1409, 13'sd2142}, {11'sd-599, 12'sd1269, 12'sd1914}},
{{12'sd2005, 13'sd-2615, 11'sd959}, {12'sd1710, 11'sd-637, 10'sd339}, {13'sd2096, 13'sd-2092, 13'sd-2635}},
{{12'sd1547, 12'sd-1478, 13'sd-2880}, {12'sd1438, 12'sd-1110, 11'sd953}, {9'sd200, 13'sd-2636, 12'sd1223}},
{{11'sd805, 13'sd2369, 13'sd-2262}, {13'sd2623, 12'sd-2030, 9'sd-173}, {12'sd-2023, 12'sd-1052, 12'sd-1294}},
{{12'sd1506, 12'sd-1982, 12'sd1287}, {11'sd785, 12'sd1757, 9'sd-233}, {12'sd1309, 11'sd-749, 12'sd1686}},
{{12'sd-1479, 13'sd2648, 12'sd1937}, {11'sd-792, 11'sd882, 12'sd-1872}, {13'sd2949, 12'sd1665, 12'sd-1867}},
{{13'sd-3141, 10'sd-367, 13'sd-2521}, {11'sd642, 13'sd-2688, 11'sd1004}, {9'sd224, 11'sd626, 12'sd-1276}}},
{
{{12'sd1281, 13'sd2100, 12'sd-1676}, {13'sd2205, 10'sd-290, 13'sd-2752}, {10'sd-448, 12'sd-1357, 10'sd351}},
{{9'sd-192, 12'sd-1309, 12'sd-1919}, {8'sd-82, 10'sd-478, 13'sd-2596}, {13'sd-2727, 11'sd912, 11'sd570}},
{{12'sd-1933, 11'sd952, 13'sd2300}, {13'sd-2357, 10'sd490, 12'sd1748}, {12'sd1238, 12'sd1736, 11'sd-993}},
{{12'sd1430, 11'sd-931, 11'sd-573}, {11'sd-722, 13'sd2552, 12'sd1913}, {12'sd1772, 12'sd1109, 9'sd-155}},
{{12'sd2010, 12'sd-1192, 12'sd1682}, {12'sd1991, 9'sd-245, 12'sd2001}, {13'sd2295, 13'sd2852, 13'sd2904}},
{{12'sd1254, 12'sd-1058, 12'sd1361}, {12'sd1394, 9'sd-132, 11'sd-667}, {12'sd1440, 12'sd1985, 13'sd-2117}},
{{13'sd3191, 12'sd1030, 12'sd-1612}, {13'sd2634, 12'sd1697, 13'sd2847}, {11'sd597, 11'sd-953, 13'sd3119}},
{{13'sd2212, 13'sd2171, 13'sd-2091}, {10'sd358, 13'sd-2390, 12'sd1361}, {12'sd1935, 12'sd-1569, 12'sd-1501}},
{{13'sd-2096, 13'sd2516, 13'sd2112}, {12'sd-1260, 12'sd1119, 12'sd-1649}, {12'sd-1165, 10'sd287, 6'sd-31}},
{{13'sd-2540, 12'sd1354, 12'sd1351}, {12'sd1294, 6'sd28, 12'sd1055}, {12'sd-1251, 13'sd2230, 13'sd2493}},
{{11'sd-705, 10'sd477, 12'sd1641}, {8'sd93, 13'sd2660, 12'sd-1155}, {11'sd-1023, 11'sd593, 12'sd1243}},
{{12'sd-1280, 12'sd1419, 10'sd424}, {11'sd957, 12'sd1103, 12'sd-1861}, {12'sd1776, 12'sd1737, 10'sd-392}},
{{7'sd54, 12'sd-2001, 11'sd-666}, {12'sd1212, 13'sd2686, 11'sd-772}, {13'sd2329, 12'sd1791, 12'sd1889}},
{{13'sd2504, 12'sd-1804, 12'sd1967}, {11'sd-1003, 12'sd-1351, 10'sd438}, {11'sd848, 12'sd1718, 8'sd-69}},
{{12'sd1308, 7'sd-43, 13'sd2184}, {13'sd2577, 13'sd3997, 12'sd1377}, {14'sd4237, 11'sd855, 13'sd2347}},
{{12'sd-1304, 11'sd942, 13'sd2211}, {12'sd-1184, 13'sd2807, 12'sd-1662}, {11'sd-655, 13'sd-2640, 13'sd2178}},
{{12'sd-1655, 13'sd2178, 12'sd1075}, {11'sd774, 11'sd-682, 11'sd-844}, {9'sd-223, 13'sd-2555, 13'sd-2536}},
{{12'sd-1389, 9'sd-193, 11'sd1021}, {12'sd1544, 12'sd-1501, 12'sd-1118}, {12'sd-1287, 11'sd-664, 10'sd-499}},
{{13'sd2635, 11'sd-573, 9'sd-238}, {13'sd2613, 7'sd57, 11'sd-862}, {11'sd-572, 13'sd2307, 13'sd-2113}},
{{12'sd1957, 12'sd1802, 13'sd-2723}, {11'sd1020, 9'sd209, 13'sd-2637}, {12'sd-1892, 13'sd-2279, 10'sd-422}},
{{13'sd2127, 10'sd472, 11'sd-524}, {10'sd402, 12'sd1848, 12'sd-1784}, {11'sd-732, 11'sd804, 10'sd257}},
{{10'sd-491, 12'sd1277, 13'sd2305}, {11'sd-712, 12'sd-1413, 12'sd-1199}, {13'sd-2269, 13'sd-2394, 12'sd-1718}},
{{9'sd220, 12'sd-1690, 8'sd92}, {13'sd2326, 7'sd46, 12'sd1112}, {11'sd-623, 13'sd2416, 11'sd992}},
{{12'sd1660, 12'sd1430, 12'sd2040}, {13'sd-2523, 13'sd2495, 11'sd848}, {12'sd-1110, 11'sd552, 12'sd-1149}},
{{12'sd1389, 11'sd-926, 11'sd725}, {12'sd-1953, 6'sd-23, 12'sd-1142}, {12'sd1919, 13'sd2086, 12'sd1953}},
{{13'sd2373, 11'sd-596, 13'sd-2245}, {12'sd-1534, 9'sd249, 12'sd1855}, {13'sd2394, 9'sd-186, 11'sd657}},
{{13'sd3306, 13'sd3379, 11'sd801}, {7'sd-36, 9'sd209, 11'sd722}, {12'sd1196, 7'sd-60, 12'sd-1425}},
{{13'sd-2200, 9'sd-245, 8'sd-72}, {13'sd2406, 12'sd1588, 12'sd-1469}, {11'sd-826, 12'sd1807, 12'sd-2044}},
{{9'sd-208, 10'sd259, 11'sd614}, {12'sd-1767, 12'sd1569, 11'sd-580}, {12'sd1979, 10'sd-452, 10'sd-386}},
{{11'sd675, 12'sd-1638, 13'sd-2859}, {10'sd-339, 12'sd-1275, 11'sd980}, {12'sd1132, 13'sd-2252, 13'sd-2656}},
{{13'sd-2349, 11'sd-531, 12'sd-1638}, {13'sd2168, 13'sd-2858, 9'sd254}, {10'sd439, 10'sd479, 11'sd-620}},
{{9'sd-166, 13'sd-2702, 12'sd1408}, {13'sd2267, 13'sd-2702, 11'sd-644}, {13'sd-2148, 13'sd-2274, 10'sd282}},
{{12'sd1115, 8'sd-112, 13'sd2694}, {12'sd-1653, 12'sd-1907, 8'sd112}, {11'sd-804, 12'sd1243, 10'sd424}},
{{12'sd1888, 12'sd1091, 9'sd163}, {13'sd-2393, 12'sd-1693, 11'sd761}, {13'sd-2503, 12'sd1742, 12'sd1701}},
{{8'sd88, 12'sd1434, 12'sd1844}, {11'sd-577, 13'sd-3202, 10'sd-372}, {12'sd1180, 10'sd289, 12'sd-1142}},
{{12'sd1555, 8'sd-85, 8'sd79}, {12'sd1170, 12'sd-1670, 10'sd-388}, {10'sd-452, 12'sd1886, 13'sd2118}},
{{12'sd-1905, 12'sd1641, 13'sd-2772}, {12'sd-2039, 13'sd-3337, 12'sd1572}, {12'sd1346, 10'sd-304, 12'sd-1079}},
{{12'sd-1215, 13'sd3211, 11'sd676}, {13'sd2649, 12'sd1589, 13'sd2330}, {13'sd2808, 10'sd-423, 13'sd2418}},
{{11'sd755, 11'sd947, 10'sd-423}, {11'sd-616, 13'sd2184, 13'sd-2188}, {11'sd890, 13'sd2523, 10'sd-486}},
{{13'sd2533, 12'sd1877, 12'sd1651}, {11'sd520, 13'sd2214, 12'sd1220}, {13'sd2459, 9'sd-222, 12'sd1867}},
{{13'sd2846, 11'sd-521, 11'sd658}, {13'sd2578, 12'sd-1433, 12'sd-1435}, {12'sd1123, 12'sd1950, 11'sd-898}},
{{12'sd1312, 13'sd-2322, 12'sd-1324}, {12'sd-1961, 12'sd1596, 9'sd217}, {12'sd-1263, 8'sd-67, 10'sd-462}},
{{13'sd2082, 13'sd2947, 12'sd-1628}, {10'sd413, 11'sd-681, 10'sd-447}, {13'sd2918, 13'sd2208, 12'sd1387}},
{{11'sd969, 12'sd-1631, 10'sd-312}, {13'sd2166, 13'sd2696, 12'sd-1535}, {12'sd1804, 13'sd3096, 12'sd1663}},
{{11'sd999, 13'sd-2678, 12'sd1475}, {11'sd1001, 10'sd-303, 13'sd-2664}, {13'sd2572, 12'sd-1975, 12'sd1509}},
{{12'sd1204, 12'sd1735, 12'sd-1727}, {13'sd-2222, 12'sd-1075, 10'sd-481}, {12'sd-1303, 13'sd-2107, 12'sd-1720}},
{{13'sd-2540, 12'sd-1511, 12'sd-1764}, {12'sd1123, 12'sd-1143, 13'sd2772}, {13'sd-2104, 13'sd-2246, 12'sd1290}},
{{10'sd365, 12'sd1041, 10'sd-387}, {11'sd-1014, 10'sd392, 12'sd1460}, {11'sd989, 11'sd763, 11'sd-756}},
{{13'sd2317, 8'sd-64, 12'sd-1588}, {12'sd1751, 10'sd450, 12'sd1673}, {12'sd-1054, 13'sd-2440, 11'sd-833}},
{{13'sd-3316, 12'sd-1126, 10'sd455}, {9'sd168, 13'sd-2415, 12'sd-1698}, {13'sd-2342, 12'sd-1333, 13'sd-2258}},
{{13'sd-2564, 12'sd-1431, 11'sd-933}, {11'sd-714, 7'sd-59, 13'sd2692}, {11'sd-929, 11'sd-533, 12'sd-1036}},
{{11'sd596, 10'sd-407, 12'sd-1390}, {13'sd-2961, 7'sd-37, 12'sd-1647}, {13'sd2497, 12'sd-1611, 7'sd49}},
{{12'sd1795, 11'sd791, 9'sd-222}, {12'sd-1498, 12'sd1179, 12'sd-1336}, {11'sd-832, 12'sd-1790, 11'sd788}},
{{11'sd850, 13'sd-2169, 12'sd-1945}, {12'sd-1726, 13'sd2673, 11'sd-755}, {9'sd-176, 10'sd-401, 13'sd2085}},
{{12'sd1284, 12'sd2034, 5'sd-10}, {12'sd-1344, 10'sd499, 12'sd1999}, {11'sd910, 13'sd2666, 12'sd-1329}},
{{13'sd-2648, 12'sd1519, 8'sd-112}, {6'sd-27, 13'sd-2688, 13'sd-2669}, {12'sd-1828, 12'sd-1936, 11'sd-650}},
{{8'sd-116, 13'sd2864, 11'sd-559}, {11'sd-792, 12'sd1424, 12'sd-1045}, {11'sd987, 14'sd4867, 12'sd1947}},
{{11'sd673, 11'sd-684, 13'sd-2261}, {11'sd-957, 13'sd-2166, 12'sd-1844}, {9'sd-248, 11'sd1005, 13'sd-2117}},
{{11'sd-830, 12'sd-1751, 13'sd2658}, {12'sd1286, 13'sd2797, 12'sd-1327}, {13'sd-2486, 10'sd381, 10'sd-369}},
{{12'sd1779, 9'sd133, 10'sd-385}, {12'sd1479, 12'sd-1435, 9'sd133}, {11'sd-977, 11'sd708, 11'sd964}},
{{7'sd-44, 12'sd1419, 12'sd-1373}, {13'sd2239, 11'sd717, 12'sd-1077}, {11'sd-1001, 13'sd-2641, 13'sd-2506}},
{{13'sd2140, 13'sd-2217, 12'sd1150}, {12'sd-1900, 13'sd-2637, 9'sd151}, {11'sd-548, 12'sd1904, 12'sd-1134}},
{{11'sd833, 12'sd-1393, 13'sd-2465}, {11'sd516, 13'sd-2487, 12'sd1460}, {12'sd1087, 9'sd-190, 13'sd2488}},
{{12'sd-1293, 12'sd1915, 11'sd591}, {13'sd-2124, 11'sd-846, 13'sd-2427}, {12'sd-1874, 9'sd135, 11'sd-601}}},
{
{{13'sd2311, 12'sd1794, 13'sd2429}, {12'sd1738, 6'sd-26, 6'sd21}, {13'sd-2065, 12'sd-1216, 11'sd-561}},
{{13'sd-2368, 12'sd-1403, 13'sd-2373}, {11'sd927, 13'sd2212, 13'sd2630}, {12'sd1519, 13'sd2592, 12'sd-1947}},
{{13'sd-2239, 4'sd4, 11'sd980}, {13'sd-2525, 13'sd-2354, 12'sd-1662}, {9'sd-133, 13'sd2539, 11'sd553}},
{{11'sd624, 12'sd1712, 13'sd2757}, {6'sd-31, 11'sd-1009, 13'sd2402}, {13'sd2477, 12'sd1294, 10'sd-284}},
{{12'sd-1706, 11'sd-892, 12'sd-1176}, {11'sd-683, 10'sd-503, 13'sd-2952}, {13'sd-2520, 8'sd-120, 12'sd-1595}},
{{10'sd510, 12'sd-1207, 14'sd4508}, {11'sd-721, 10'sd464, 12'sd1934}, {13'sd-3415, 11'sd-576, 13'sd3016}},
{{13'sd-2996, 11'sd-1022, 6'sd16}, {13'sd-3757, 13'sd-2667, 11'sd737}, {12'sd-1409, 8'sd-110, 8'sd74}},
{{13'sd2450, 10'sd-496, 8'sd117}, {12'sd1965, 13'sd-2421, 11'sd700}, {12'sd-1299, 12'sd-1873, 12'sd1507}},
{{12'sd1944, 9'sd-179, 13'sd-2743}, {11'sd-851, 13'sd-2485, 12'sd1222}, {6'sd19, 11'sd627, 12'sd1151}},
{{12'sd1864, 13'sd-2218, 11'sd-571}, {13'sd2467, 10'sd-279, 12'sd1202}, {13'sd2229, 12'sd1084, 7'sd43}},
{{11'sd-549, 9'sd-238, 13'sd-2451}, {10'sd363, 13'sd-3150, 12'sd1592}, {12'sd1541, 13'sd-2281, 11'sd594}},
{{10'sd359, 13'sd2272, 12'sd1540}, {13'sd-2320, 9'sd167, 13'sd2763}, {12'sd-1476, 13'sd2431, 12'sd1144}},
{{12'sd-1354, 12'sd1134, 13'sd-3025}, {12'sd-1783, 11'sd-674, 12'sd-1358}, {11'sd-987, 12'sd2031, 13'sd-2115}},
{{11'sd957, 12'sd1097, 12'sd-1506}, {13'sd2463, 12'sd1117, 12'sd-1801}, {13'sd2482, 13'sd-2843, 11'sd-819}},
{{11'sd-936, 10'sd-265, 12'sd1605}, {13'sd-2763, 9'sd-249, 11'sd779}, {13'sd-2475, 12'sd1066, 12'sd-1422}},
{{12'sd-2032, 12'sd1592, 11'sd896}, {12'sd1384, 4'sd-6, 8'sd-67}, {13'sd-2626, 12'sd-1848, 12'sd-1721}},
{{11'sd665, 12'sd-1961, 12'sd1877}, {11'sd-904, 13'sd2566, 12'sd1371}, {13'sd2189, 13'sd-2149, 13'sd2303}},
{{12'sd-2006, 13'sd-2518, 7'sd-51}, {13'sd-3200, 12'sd1972, 13'sd-2746}, {13'sd-2097, 13'sd-2127, 5'sd-9}},
{{11'sd-741, 12'sd-1107, 12'sd1137}, {10'sd334, 11'sd791, 10'sd-284}, {12'sd-1361, 12'sd-1712, 10'sd506}},
{{12'sd1474, 13'sd2486, 12'sd-1387}, {12'sd-1344, 12'sd1069, 11'sd933}, {13'sd2156, 12'sd-1651, 11'sd-1013}},
{{12'sd1036, 9'sd167, 11'sd582}, {13'sd2433, 12'sd-1424, 12'sd-1779}, {12'sd-1879, 12'sd-1901, 13'sd-2184}},
{{13'sd3078, 13'sd2670, 7'sd37}, {13'sd2973, 12'sd-1697, 12'sd-1393}, {10'sd324, 12'sd1310, 13'sd2186}},
{{12'sd-2031, 8'sd-126, 12'sd-1388}, {12'sd1039, 12'sd-1253, 3'sd3}, {11'sd729, 9'sd-128, 12'sd-1413}},
{{10'sd301, 10'sd447, 13'sd-2090}, {13'sd2471, 12'sd-1177, 7'sd-32}, {12'sd1440, 10'sd321, 12'sd-1507}},
{{11'sd-609, 13'sd2211, 12'sd1707}, {12'sd1197, 13'sd2572, 9'sd-179}, {13'sd2253, 12'sd1164, 13'sd2451}},
{{12'sd1749, 9'sd-140, 13'sd2104}, {11'sd-543, 13'sd-2161, 12'sd-1352}, {12'sd1550, 12'sd-1966, 12'sd1127}},
{{13'sd-2393, 13'sd2224, 10'sd-386}, {12'sd1849, 13'sd3485, 12'sd-1186}, {10'sd-451, 13'sd3233, 13'sd2501}},
{{12'sd1502, 9'sd-168, 13'sd2211}, {13'sd2377, 12'sd-1528, 13'sd-2215}, {11'sd-592, 11'sd988, 11'sd797}},
{{13'sd2578, 13'sd2420, 12'sd1658}, {12'sd1118, 8'sd87, 11'sd-553}, {11'sd-920, 13'sd-2512, 12'sd1920}},
{{12'sd-1912, 10'sd-441, 8'sd86}, {11'sd-579, 11'sd906, 12'sd2027}, {13'sd-2253, 13'sd-2205, 13'sd-2343}},
{{9'sd-212, 12'sd-1334, 12'sd1805}, {9'sd163, 12'sd-1464, 7'sd-51}, {12'sd1284, 11'sd-523, 13'sd-2092}},
{{13'sd-2252, 11'sd577, 12'sd1531}, {13'sd2495, 10'sd-477, 12'sd1936}, {11'sd-989, 11'sd-532, 11'sd512}},
{{11'sd643, 12'sd-1792, 11'sd999}, {12'sd-1351, 12'sd-1250, 13'sd-2899}, {13'sd2594, 11'sd-743, 12'sd-1458}},
{{13'sd-3103, 13'sd-2340, 13'sd-2157}, {12'sd1140, 11'sd-533, 11'sd597}, {13'sd2209, 13'sd2207, 9'sd-228}},
{{12'sd1785, 12'sd1341, 10'sd382}, {11'sd530, 12'sd1622, 10'sd404}, {11'sd753, 9'sd162, 9'sd139}},
{{12'sd-1313, 12'sd1539, 12'sd1350}, {13'sd2096, 10'sd-383, 9'sd-162}, {13'sd2212, 12'sd1600, 12'sd-1201}},
{{11'sd-531, 12'sd-1434, 11'sd-1008}, {11'sd621, 11'sd-841, 12'sd1568}, {13'sd2184, 10'sd-384, 12'sd1035}},
{{12'sd-1831, 13'sd2667, 11'sd-575}, {11'sd-617, 12'sd2034, 11'sd873}, {12'sd-1602, 12'sd-1361, 13'sd2537}},
{{11'sd-570, 12'sd-1251, 12'sd1650}, {12'sd-1626, 12'sd-1939, 11'sd554}, {13'sd2993, 13'sd2797, 13'sd2310}},
{{13'sd-2496, 13'sd2083, 13'sd2264}, {12'sd-1729, 7'sd-37, 12'sd-1831}, {13'sd2390, 11'sd629, 12'sd2031}},
{{9'sd-134, 11'sd-756, 11'sd-767}, {11'sd566, 11'sd934, 8'sd-66}, {10'sd-351, 11'sd845, 12'sd-1934}},
{{12'sd-1127, 13'sd2907, 13'sd2121}, {12'sd-1095, 13'sd-2428, 11'sd522}, {12'sd1830, 11'sd749, 13'sd-2256}},
{{11'sd710, 11'sd-683, 12'sd1769}, {12'sd1835, 11'sd-681, 12'sd-1756}, {12'sd1167, 11'sd-1004, 13'sd-2453}},
{{11'sd936, 12'sd1160, 11'sd957}, {12'sd1659, 12'sd1651, 13'sd3886}, {13'sd3059, 12'sd1419, 12'sd1082}},
{{12'sd1896, 12'sd1177, 10'sd505}, {11'sd-997, 9'sd-132, 13'sd2234}, {13'sd-2484, 13'sd-2081, 13'sd2630}},
{{13'sd2342, 12'sd1909, 11'sd-832}, {8'sd-102, 10'sd274, 10'sd-342}, {12'sd1091, 12'sd1347, 13'sd2473}},
{{12'sd-1623, 12'sd-1509, 6'sd24}, {13'sd-2640, 10'sd-272, 12'sd1623}, {13'sd2528, 13'sd3016, 11'sd542}},
{{10'sd316, 13'sd-2132, 12'sd1493}, {12'sd1739, 13'sd-2514, 11'sd-731}, {9'sd239, 12'sd-1865, 13'sd-2406}},
{{10'sd478, 10'sd-258, 12'sd-1849}, {13'sd2075, 13'sd2188, 13'sd2110}, {13'sd-2148, 10'sd453, 12'sd1887}},
{{13'sd2215, 12'sd-1275, 12'sd-1882}, {12'sd1675, 10'sd-317, 11'sd-1008}, {13'sd-2997, 9'sd-221, 8'sd-105}},
{{11'sd-988, 12'sd-1407, 13'sd-2242}, {12'sd-1181, 13'sd-2129, 11'sd666}, {13'sd-2050, 10'sd-311, 13'sd-2553}},
{{13'sd2710, 12'sd-1882, 12'sd-1701}, {12'sd1143, 12'sd1860, 9'sd241}, {12'sd-1539, 11'sd531, 13'sd2213}},
{{12'sd1213, 12'sd1044, 13'sd-2351}, {12'sd1236, 13'sd-2538, 12'sd-1715}, {12'sd1543, 13'sd-2667, 12'sd-1551}},
{{8'sd110, 12'sd1902, 11'sd948}, {8'sd96, 11'sd-798, 11'sd-800}, {12'sd-1042, 12'sd-1214, 12'sd-1039}},
{{12'sd1585, 12'sd1452, 11'sd855}, {12'sd-1834, 11'sd-860, 13'sd-2613}, {10'sd467, 11'sd793, 13'sd-2127}},
{{12'sd-1796, 13'sd2420, 11'sd720}, {12'sd1753, 12'sd1400, 10'sd-404}, {13'sd-2255, 12'sd1829, 12'sd-1333}},
{{10'sd292, 10'sd472, 12'sd1456}, {11'sd-914, 13'sd-2605, 13'sd-2263}, {12'sd-1329, 11'sd-624, 11'sd-793}},
{{12'sd-1520, 10'sd418, 13'sd2094}, {10'sd300, 12'sd-1385, 13'sd-2132}, {11'sd-910, 13'sd2309, 11'sd625}},
{{12'sd2019, 13'sd-2661, 12'sd-1698}, {13'sd2065, 12'sd1964, 13'sd-2050}, {12'sd1645, 12'sd1964, 13'sd2240}},
{{13'sd-2533, 11'sd-979, 13'sd3420}, {8'sd65, 12'sd-1855, 10'sd-309}, {13'sd-2171, 13'sd-2105, 13'sd2669}},
{{11'sd-570, 10'sd293, 10'sd293}, {12'sd-1435, 12'sd1643, 11'sd622}, {13'sd-2105, 11'sd-858, 9'sd-179}},
{{13'sd2871, 13'sd2303, 9'sd210}, {12'sd1836, 9'sd132, 12'sd-1026}, {13'sd-2122, 11'sd-1001, 12'sd-1551}},
{{11'sd863, 12'sd1727, 11'sd879}, {12'sd-1304, 11'sd-706, 13'sd2242}, {11'sd-932, 13'sd2930, 6'sd25}},
{{11'sd976, 13'sd2091, 11'sd610}, {11'sd981, 12'sd-1139, 11'sd-526}, {12'sd-1251, 11'sd773, 12'sd1712}}},
{
{{13'sd2618, 12'sd-1177, 7'sd52}, {9'sd-199, 11'sd711, 13'sd-2439}, {12'sd1086, 11'sd517, 12'sd-1658}},
{{13'sd2700, 12'sd1091, 10'sd403}, {12'sd1374, 12'sd-1280, 8'sd-92}, {14'sd4140, 10'sd-416, 13'sd3239}},
{{13'sd-2683, 11'sd-951, 10'sd-435}, {12'sd-1845, 13'sd2366, 12'sd2022}, {11'sd-566, 12'sd1577, 12'sd1849}},
{{13'sd-2148, 11'sd679, 13'sd2386}, {12'sd-1459, 5'sd-11, 13'sd2218}, {11'sd947, 11'sd856, 12'sd-1440}},
{{13'sd2480, 11'sd-644, 13'sd3503}, {11'sd-556, 11'sd702, 13'sd3031}, {13'sd-2365, 12'sd-1182, 11'sd910}},
{{11'sd739, 13'sd2382, 13'sd3223}, {10'sd-379, 8'sd85, 14'sd4286}, {11'sd-669, 13'sd2911, 11'sd-672}},
{{13'sd-2841, 11'sd1007, 13'sd2246}, {14'sd-4744, 12'sd-1345, 12'sd1898}, {14'sd-4243, 11'sd-541, 13'sd4059}},
{{12'sd-1055, 12'sd-1252, 13'sd2666}, {12'sd-1225, 13'sd2528, 13'sd3211}, {13'sd-2320, 9'sd241, 10'sd429}},
{{11'sd694, 12'sd-1687, 8'sd-125}, {12'sd1464, 13'sd2485, 11'sd820}, {12'sd-2040, 12'sd-1846, 13'sd-2535}},
{{11'sd972, 11'sd-801, 12'sd1986}, {13'sd2373, 11'sd-519, 11'sd-844}, {11'sd1022, 11'sd-863, 8'sd-105}},
{{9'sd-228, 13'sd-2999, 13'sd2065}, {13'sd-2561, 12'sd1323, 12'sd1978}, {12'sd-1779, 12'sd-1878, 11'sd881}},
{{13'sd2216, 11'sd918, 10'sd279}, {10'sd271, 10'sd451, 13'sd-2271}, {11'sd807, 10'sd379, 12'sd1885}},
{{12'sd1027, 13'sd3188, 12'sd1851}, {13'sd2758, 10'sd-302, 8'sd-121}, {13'sd3582, 13'sd3536, 12'sd1229}},
{{12'sd1145, 12'sd-2015, 12'sd1362}, {12'sd-1657, 13'sd2449, 12'sd1418}, {12'sd-1031, 11'sd589, 11'sd932}},
{{13'sd-2236, 14'sd-6147, 11'sd-1017}, {14'sd-5431, 13'sd-3185, 13'sd-2361}, {15'sd-9563, 14'sd-6413, 13'sd-4017}},
{{11'sd542, 12'sd1465, 13'sd-2541}, {9'sd185, 11'sd-1013, 12'sd1549}, {14'sd4597, 11'sd-734, 12'sd1253}},
{{12'sd1309, 13'sd2058, 13'sd-2210}, {12'sd-1222, 11'sd767, 12'sd1154}, {12'sd-1193, 12'sd-1648, 12'sd-1593}},
{{11'sd-889, 10'sd-463, 12'sd1551}, {12'sd1909, 11'sd-991, 13'sd3268}, {13'sd-3183, 11'sd1008, 13'sd3642}},
{{12'sd1706, 11'sd781, 13'sd-2735}, {11'sd1021, 12'sd-1249, 12'sd1121}, {12'sd-1478, 13'sd2335, 13'sd2295}},
{{10'sd-457, 12'sd1129, 6'sd19}, {12'sd1269, 12'sd-2032, 10'sd-284}, {12'sd-1970, 12'sd1269, 13'sd-3155}},
{{11'sd761, 10'sd292, 12'sd1903}, {12'sd1591, 12'sd1697, 13'sd-2885}, {10'sd316, 12'sd-1238, 13'sd-2837}},
{{11'sd993, 10'sd-397, 12'sd1175}, {11'sd1018, 12'sd-1530, 11'sd-766}, {12'sd1911, 13'sd2766, 13'sd-2500}},
{{12'sd1436, 12'sd-1513, 10'sd437}, {13'sd2624, 13'sd2939, 13'sd2682}, {13'sd2390, 12'sd1361, 13'sd3041}},
{{13'sd-3164, 11'sd-677, 12'sd-1608}, {8'sd-79, 10'sd-278, 13'sd-2953}, {13'sd-2424, 12'sd1053, 12'sd-1127}},
{{12'sd-1647, 12'sd1543, 12'sd1290}, {11'sd-940, 12'sd1978, 11'sd695}, {13'sd2635, 13'sd-2081, 11'sd-966}},
{{12'sd1060, 11'sd736, 12'sd-1804}, {11'sd975, 12'sd1839, 13'sd2340}, {13'sd2695, 13'sd-2153, 13'sd2316}},
{{14'sd-5330, 13'sd-2933, 13'sd2431}, {13'sd-3940, 8'sd-77, 11'sd762}, {14'sd-4099, 12'sd1964, 8'sd89}},
{{12'sd-1090, 11'sd517, 12'sd1989}, {12'sd1473, 13'sd-2545, 13'sd-3523}, {10'sd-508, 13'sd-4011, 13'sd-3271}},
{{12'sd-1829, 13'sd-2412, 13'sd-2337}, {13'sd-2983, 12'sd-1605, 11'sd905}, {12'sd-1784, 13'sd-3684, 11'sd-813}},
{{11'sd628, 13'sd-2980, 9'sd240}, {10'sd-417, 11'sd-791, 13'sd-2724}, {11'sd765, 11'sd1019, 12'sd1818}},
{{12'sd1952, 13'sd2538, 12'sd-1129}, {10'sd445, 11'sd-707, 12'sd-1164}, {12'sd-1953, 10'sd-473, 13'sd2534}},
{{13'sd3029, 12'sd-1081, 12'sd-1502}, {13'sd3165, 12'sd1952, 12'sd1530}, {12'sd-1643, 11'sd-851, 12'sd-1080}},
{{12'sd1771, 9'sd169, 12'sd1991}, {11'sd685, 11'sd-985, 13'sd-2934}, {12'sd1589, 10'sd-464, 13'sd-2630}},
{{11'sd-603, 13'sd-2230, 13'sd-3559}, {12'sd1038, 11'sd-746, 12'sd-1418}, {13'sd-2627, 12'sd-2009, 11'sd-1012}},
{{10'sd272, 13'sd-2417, 11'sd-517}, {12'sd1173, 11'sd579, 13'sd-3428}, {11'sd-623, 12'sd2027, 13'sd-2532}},
{{12'sd-1278, 13'sd2705, 13'sd-2359}, {11'sd947, 13'sd2557, 13'sd-2508}, {13'sd2295, 12'sd1608, 11'sd-631}},
{{11'sd-975, 12'sd-1656, 12'sd-1643}, {12'sd-1983, 13'sd-4067, 13'sd-2865}, {13'sd-2659, 9'sd225, 12'sd-1857}},
{{12'sd-1154, 13'sd3549, 13'sd2196}, {13'sd-3408, 9'sd172, 13'sd2338}, {12'sd1476, 13'sd3117, 13'sd3981}},
{{13'sd-2924, 11'sd-661, 13'sd2842}, {10'sd364, 11'sd-582, 13'sd2706}, {10'sd348, 10'sd-312, 13'sd2503}},
{{12'sd-1386, 12'sd1655, 12'sd1675}, {12'sd1518, 10'sd256, 10'sd-511}, {10'sd300, 12'sd1974, 12'sd1956}},
{{13'sd-2745, 11'sd-905, 11'sd-656}, {13'sd-2376, 11'sd-1021, 12'sd1625}, {12'sd-1987, 12'sd-1212, 13'sd2243}},
{{13'sd2381, 10'sd-431, 12'sd2003}, {11'sd974, 11'sd652, 13'sd2306}, {12'sd1950, 12'sd-1080, 12'sd1593}},
{{12'sd-1318, 14'sd-4513, 13'sd2727}, {14'sd-6639, 13'sd-2637, 13'sd-2598}, {14'sd-5231, 11'sd-725, 7'sd-56}},
{{12'sd-1087, 11'sd705, 14'sd5011}, {10'sd-338, 14'sd4918, 13'sd2654}, {13'sd2604, 14'sd6692, 14'sd5209}},
{{10'sd-330, 11'sd969, 12'sd-1552}, {12'sd-1979, 10'sd-263, 12'sd1395}, {11'sd1011, 12'sd-1313, 12'sd1331}},
{{12'sd-1935, 11'sd-718, 11'sd-953}, {13'sd2160, 13'sd3123, 11'sd806}, {13'sd2864, 13'sd3130, 12'sd-1490}},
{{11'sd702, 12'sd-1544, 13'sd-4049}, {13'sd2198, 11'sd927, 12'sd-1998}, {11'sd-956, 11'sd625, 13'sd-2806}},
{{13'sd-3037, 13'sd-2819, 8'sd-127}, {10'sd-327, 13'sd-3451, 12'sd2031}, {12'sd-1178, 12'sd-1770, 10'sd-336}},
{{13'sd-3792, 12'sd1308, 13'sd-2590}, {9'sd192, 14'sd-4151, 11'sd-875}, {8'sd-76, 13'sd-2334, 13'sd2171}},
{{13'sd2949, 13'sd-2266, 12'sd-2035}, {14'sd4622, 12'sd1328, 12'sd-1627}, {12'sd1264, 13'sd2709, 9'sd185}},
{{11'sd574, 12'sd1583, 12'sd-1364}, {13'sd2065, 12'sd1182, 12'sd1849}, {13'sd-2235, 13'sd-2561, 12'sd1144}},
{{12'sd-1987, 7'sd-39, 9'sd232}, {12'sd-1951, 11'sd773, 13'sd-2410}, {11'sd-626, 12'sd-1286, 11'sd-971}},
{{9'sd-182, 13'sd2138, 13'sd-2739}, {13'sd-2934, 13'sd-2274, 12'sd1981}, {13'sd-2718, 13'sd-2174, 11'sd-936}},
{{10'sd-390, 12'sd-1971, 13'sd2222}, {12'sd-1717, 7'sd-51, 9'sd-253}, {13'sd2329, 13'sd2753, 12'sd1206}},
{{11'sd-929, 13'sd-2441, 6'sd18}, {13'sd-2605, 11'sd536, 12'sd1910}, {13'sd-3004, 12'sd2006, 12'sd1456}},
{{13'sd-2703, 6'sd31, 12'sd-1036}, {13'sd-2435, 11'sd-992, 12'sd1388}, {12'sd1814, 12'sd-1182, 11'sd-909}},
{{11'sd988, 11'sd514, 13'sd2354}, {10'sd393, 12'sd1900, 13'sd2187}, {12'sd-1537, 12'sd1145, 12'sd-1351}},
{{13'sd2766, 12'sd-1269, 12'sd-1331}, {8'sd-113, 12'sd-1419, 13'sd2526}, {11'sd571, 11'sd650, 13'sd3008}},
{{12'sd1450, 10'sd-342, 13'sd2061}, {13'sd-2279, 11'sd-613, 11'sd903}, {10'sd-424, 11'sd-782, 11'sd-818}},
{{12'sd1583, 13'sd-2081, 10'sd327}, {14'sd-5225, 13'sd-3793, 11'sd-866}, {12'sd-1618, 11'sd-791, 13'sd-2689}},
{{13'sd2522, 11'sd571, 13'sd-2503}, {13'sd2858, 11'sd953, 12'sd1841}, {11'sd607, 11'sd729, 11'sd-686}},
{{13'sd3445, 12'sd-1581, 13'sd-2698}, {5'sd-9, 9'sd154, 12'sd-1389}, {13'sd-2077, 7'sd-47, 13'sd-2672}},
{{13'sd2205, 12'sd-1612, 12'sd1244}, {13'sd2269, 12'sd1330, 13'sd2264}, {11'sd-622, 11'sd-564, 11'sd-895}},
{{10'sd-418, 9'sd203, 12'sd-1863}, {13'sd-2657, 14'sd-4208, 12'sd1109}, {13'sd-2300, 8'sd68, 12'sd1170}}},
{
{{12'sd-1150, 8'sd-97, 13'sd2274}, {12'sd1526, 12'sd1381, 13'sd2513}, {12'sd-1248, 13'sd-2413, 13'sd-2349}},
{{13'sd-2505, 12'sd1087, 12'sd1760}, {12'sd-1256, 12'sd-1255, 13'sd2808}, {13'sd2863, 12'sd-1548, 11'sd996}},
{{12'sd-1234, 13'sd-2937, 12'sd-1234}, {13'sd-2330, 9'sd-177, 13'sd2624}, {11'sd-547, 8'sd121, 12'sd1245}},
{{12'sd-1456, 13'sd-2945, 10'sd-284}, {12'sd-1806, 13'sd-2344, 12'sd1573}, {9'sd177, 12'sd1141, 11'sd850}},
{{11'sd-554, 13'sd2850, 13'sd3330}, {11'sd-616, 14'sd4540, 10'sd492}, {13'sd-2203, 8'sd-76, 11'sd532}},
{{9'sd-234, 13'sd3379, 11'sd602}, {12'sd-1510, 10'sd355, 12'sd1460}, {10'sd-423, 13'sd2692, 12'sd1136}},
{{9'sd-195, 12'sd1900, 13'sd2137}, {11'sd-586, 10'sd-497, 13'sd-3775}, {12'sd-1277, 11'sd895, 13'sd-3779}},
{{12'sd-1378, 13'sd2290, 11'sd705}, {7'sd59, 13'sd-2862, 12'sd2018}, {9'sd252, 11'sd-986, 12'sd-1611}},
{{11'sd536, 13'sd2627, 11'sd-744}, {10'sd-264, 11'sd-790, 10'sd265}, {13'sd2071, 10'sd497, 10'sd381}},
{{12'sd-1268, 11'sd782, 12'sd1048}, {10'sd507, 12'sd-1808, 6'sd30}, {13'sd-3166, 12'sd-1575, 13'sd-2582}},
{{12'sd1284, 11'sd-843, 12'sd1135}, {12'sd-1065, 13'sd-2255, 11'sd-809}, {12'sd-1987, 9'sd-189, 12'sd-1238}},
{{9'sd-166, 13'sd-2822, 11'sd-545}, {12'sd1468, 12'sd-1654, 10'sd-371}, {10'sd-469, 12'sd-1256, 12'sd-1551}},
{{13'sd3033, 11'sd602, 9'sd224}, {12'sd-1112, 8'sd-124, 10'sd375}, {12'sd1362, 10'sd477, 13'sd3021}},
{{13'sd2728, 13'sd-3143, 13'sd-3151}, {12'sd1742, 12'sd-1837, 13'sd-2473}, {11'sd-575, 12'sd-1876, 12'sd-1949}},
{{3'sd-3, 11'sd905, 11'sd-998}, {13'sd-3492, 8'sd-94, 13'sd-3104}, {13'sd-2543, 14'sd-5751, 14'sd-5276}},
{{8'sd115, 12'sd-1068, 12'sd1368}, {11'sd715, 11'sd-556, 11'sd-614}, {13'sd3662, 12'sd-1243, 14'sd4256}},
{{13'sd2238, 10'sd-431, 11'sd519}, {13'sd2590, 13'sd2141, 13'sd-2433}, {11'sd963, 12'sd1899, 13'sd-2362}},
{{13'sd2773, 12'sd-1189, 13'sd2888}, {12'sd1144, 12'sd-1480, 13'sd3708}, {12'sd1347, 9'sd-160, 11'sd-527}},
{{13'sd2559, 10'sd433, 13'sd-2224}, {12'sd1979, 12'sd1242, 13'sd-2581}, {12'sd1684, 13'sd-2660, 13'sd-2538}},
{{12'sd1854, 13'sd-2627, 13'sd-2914}, {12'sd1773, 9'sd-218, 10'sd-273}, {10'sd-276, 10'sd-276, 12'sd-1723}},
{{12'sd1451, 12'sd-1432, 12'sd-1223}, {13'sd2663, 9'sd208, 13'sd-3083}, {12'sd1487, 13'sd-2229, 12'sd-1979}},
{{12'sd-1159, 13'sd2228, 12'sd1232}, {13'sd2781, 11'sd-602, 12'sd1371}, {10'sd422, 12'sd-1029, 12'sd-1235}},
{{12'sd-1463, 7'sd42, 13'sd2064}, {13'sd3020, 12'sd2014, 12'sd-1266}, {13'sd2765, 13'sd2243, 12'sd-1550}},
{{13'sd-2222, 13'sd-2102, 11'sd-762}, {12'sd1208, 13'sd2152, 12'sd-1287}, {13'sd-2353, 12'sd-1693, 11'sd593}},
{{10'sd412, 12'sd-1375, 12'sd1204}, {11'sd-992, 13'sd2436, 11'sd726}, {9'sd-136, 12'sd1344, 12'sd1845}},
{{8'sd108, 11'sd855, 12'sd1960}, {2'sd-1, 12'sd1802, 11'sd-653}, {13'sd2072, 10'sd407, 10'sd-370}},
{{11'sd618, 13'sd-3216, 7'sd-36}, {11'sd601, 10'sd278, 11'sd594}, {14'sd4554, 13'sd2048, 12'sd-1667}},
{{11'sd989, 12'sd1406, 12'sd-1041}, {11'sd-784, 12'sd-1305, 5'sd15}, {13'sd-2302, 11'sd856, 13'sd-2417}},
{{10'sd265, 3'sd3, 12'sd-1774}, {13'sd-2768, 13'sd-2665, 11'sd699}, {12'sd-1589, 11'sd-898, 9'sd-165}},
{{12'sd-1187, 12'sd-1659, 11'sd-517}, {12'sd-1568, 12'sd1321, 12'sd-1294}, {13'sd2198, 11'sd708, 12'sd2035}},
{{8'sd-65, 12'sd1618, 11'sd-941}, {12'sd1820, 12'sd-1917, 12'sd-1467}, {13'sd2351, 12'sd-1785, 12'sd-1290}},
{{12'sd1138, 12'sd-1223, 13'sd-2150}, {10'sd289, 12'sd1390, 11'sd-691}, {13'sd2317, 13'sd-2064, 11'sd-871}},
{{12'sd-1066, 12'sd1728, 11'sd-816}, {12'sd1558, 13'sd2115, 8'sd106}, {12'sd1464, 12'sd-1632, 11'sd-536}},
{{11'sd648, 9'sd238, 11'sd-988}, {13'sd-2674, 11'sd-966, 11'sd928}, {11'sd870, 12'sd1391, 13'sd-2817}},
{{10'sd-344, 12'sd1358, 10'sd-399}, {10'sd443, 12'sd1116, 11'sd551}, {12'sd1267, 11'sd-748, 11'sd611}},
{{9'sd200, 11'sd942, 11'sd821}, {12'sd2036, 12'sd-1317, 12'sd-1105}, {10'sd-482, 12'sd1343, 11'sd-976}},
{{12'sd-1631, 13'sd2049, 10'sd464}, {11'sd851, 11'sd838, 13'sd-3656}, {13'sd2671, 13'sd2214, 13'sd-2791}},
{{12'sd-1623, 9'sd165, 12'sd-1181}, {12'sd1603, 12'sd-1759, 11'sd-911}, {13'sd3650, 13'sd3411, 8'sd113}},
{{8'sd93, 12'sd-1908, 12'sd-1270}, {13'sd2424, 12'sd-1249, 13'sd-2370}, {13'sd-2201, 8'sd-93, 12'sd1104}},
{{12'sd-1390, 11'sd-860, 12'sd-1043}, {13'sd2486, 13'sd2769, 9'sd-131}, {13'sd-2676, 11'sd-840, 12'sd1035}},
{{12'sd1672, 13'sd3278, 12'sd1393}, {13'sd2482, 12'sd-1643, 10'sd260}, {13'sd3168, 13'sd2772, 11'sd744}},
{{12'sd1553, 11'sd-818, 12'sd1434}, {12'sd-1332, 12'sd1946, 11'sd-651}, {12'sd-2009, 13'sd2065, 10'sd360}},
{{12'sd-1703, 13'sd-2849, 11'sd735}, {10'sd-298, 13'sd-3438, 13'sd-2563}, {12'sd-1804, 13'sd-3960, 13'sd-3385}},
{{13'sd-3321, 12'sd-1768, 13'sd-3204}, {13'sd4094, 12'sd1267, 12'sd-1678}, {14'sd7513, 13'sd3736, 13'sd3494}},
{{11'sd-882, 8'sd99, 12'sd1525}, {12'sd1976, 11'sd649, 13'sd2372}, {12'sd1394, 12'sd1545, 11'sd-563}},
{{12'sd-1319, 13'sd2139, 12'sd1407}, {8'sd-93, 12'sd1319, 11'sd587}, {12'sd1341, 11'sd-515, 13'sd2351}},
{{12'sd1978, 12'sd1582, 12'sd-1473}, {11'sd735, 11'sd1019, 10'sd-504}, {14'sd4386, 11'sd-950, 13'sd2965}},
{{13'sd2465, 13'sd-2545, 13'sd-3168}, {13'sd2819, 12'sd-1387, 12'sd1071}, {12'sd1601, 12'sd-1111, 11'sd758}},
{{10'sd-455, 12'sd-1441, 13'sd-3117}, {12'sd-1739, 13'sd-2265, 13'sd-2306}, {13'sd-2527, 10'sd425, 10'sd294}},
{{8'sd91, 9'sd-232, 10'sd390}, {7'sd-40, 13'sd3465, 13'sd2779}, {8'sd91, 9'sd252, 11'sd-985}},
{{13'sd-2124, 12'sd1302, 13'sd-2841}, {13'sd2234, 12'sd-1219, 12'sd1558}, {12'sd1113, 12'sd-1828, 13'sd2528}},
{{11'sd-568, 13'sd-2502, 13'sd2473}, {12'sd1555, 6'sd23, 12'sd-1566}, {12'sd-1937, 9'sd190, 11'sd804}},
{{11'sd-936, 12'sd1861, 11'sd550}, {12'sd1202, 11'sd521, 12'sd1313}, {13'sd-2474, 14'sd-5879, 13'sd-3828}},
{{11'sd649, 12'sd-1434, 7'sd62}, {10'sd325, 13'sd-2728, 13'sd-2846}, {11'sd587, 5'sd-13, 6'sd18}},
{{11'sd847, 13'sd3085, 14'sd4872}, {11'sd882, 12'sd2012, 13'sd3924}, {12'sd-1037, 12'sd-1225, 11'sd979}},
{{12'sd-1301, 13'sd2327, 13'sd-2873}, {13'sd2109, 11'sd785, 11'sd-968}, {10'sd-360, 13'sd-2454, 11'sd759}},
{{11'sd958, 13'sd-2059, 14'sd4193}, {12'sd-1943, 12'sd-1661, 13'sd3031}, {13'sd-3486, 14'sd-5160, 12'sd1038}},
{{10'sd-382, 12'sd-1576, 5'sd-13}, {12'sd1800, 13'sd3380, 10'sd407}, {11'sd-992, 13'sd2430, 8'sd-84}},
{{13'sd-2715, 12'sd1583, 11'sd584}, {10'sd-404, 12'sd1125, 9'sd251}, {12'sd1704, 13'sd-2711, 11'sd537}},
{{13'sd2253, 12'sd1367, 12'sd1667}, {12'sd1146, 11'sd837, 10'sd-299}, {13'sd2175, 12'sd1027, 12'sd1872}},
{{10'sd509, 12'sd1973, 12'sd-1728}, {9'sd-130, 11'sd777, 10'sd342}, {10'sd-362, 12'sd1920, 12'sd-1460}},
{{12'sd1277, 12'sd1804, 12'sd-1211}, {12'sd-1240, 11'sd801, 12'sd1731}, {12'sd-1298, 10'sd262, 12'sd-1969}},
{{11'sd656, 12'sd1976, 10'sd358}, {10'sd-369, 11'sd-913, 12'sd-1823}, {13'sd3233, 11'sd-918, 9'sd-238}},
{{14'sd-4240, 14'sd-4375, 14'sd-4366}, {13'sd-3240, 13'sd-2698, 14'sd-4735}, {14'sd-4248, 14'sd-4365, 12'sd-1389}}},
{
{{13'sd-2117, 13'sd2420, 11'sd-538}, {13'sd-3181, 10'sd-395, 12'sd-1594}, {11'sd816, 13'sd2064, 8'sd90}},
{{10'sd292, 12'sd-1590, 11'sd971}, {11'sd-978, 11'sd718, 12'sd-1640}, {12'sd1411, 12'sd-2022, 12'sd1409}},
{{11'sd885, 13'sd2633, 11'sd965}, {13'sd2077, 12'sd1245, 11'sd747}, {13'sd2291, 13'sd-2692, 13'sd2224}},
{{13'sd2159, 12'sd-1751, 8'sd-120}, {12'sd1198, 12'sd2035, 10'sd355}, {12'sd1972, 13'sd-2625, 12'sd-1967}},
{{14'sd6797, 14'sd5792, 10'sd-426}, {13'sd3980, 11'sd616, 11'sd951}, {13'sd-2404, 11'sd907, 12'sd1182}},
{{13'sd3062, 12'sd1259, 10'sd-489}, {13'sd-3468, 11'sd-522, 12'sd1202}, {10'sd412, 12'sd-1372, 13'sd2106}},
{{12'sd-1160, 13'sd-2999, 13'sd-3039}, {13'sd-2892, 10'sd-437, 11'sd-925}, {11'sd-986, 10'sd343, 9'sd237}},
{{10'sd261, 12'sd-1943, 11'sd709}, {13'sd-2449, 13'sd-2404, 11'sd514}, {13'sd2418, 12'sd-1605, 11'sd720}},
{{12'sd1075, 12'sd-1292, 12'sd-1883}, {12'sd1153, 13'sd-2682, 11'sd-1002}, {12'sd-1648, 11'sd-986, 12'sd1526}},
{{13'sd-2075, 13'sd-2320, 7'sd-39}, {13'sd-2290, 12'sd1792, 11'sd-693}, {10'sd-384, 11'sd667, 10'sd-457}},
{{12'sd-1686, 12'sd-1769, 11'sd1010}, {12'sd-1724, 8'sd125, 10'sd434}, {12'sd-1442, 5'sd-13, 11'sd-562}},
{{12'sd1407, 13'sd2897, 13'sd2512}, {10'sd-336, 12'sd-1219, 12'sd1033}, {11'sd621, 11'sd987, 12'sd1563}},
{{9'sd153, 13'sd2083, 13'sd-2332}, {12'sd-1637, 13'sd-2561, 11'sd-858}, {13'sd2113, 11'sd889, 12'sd-1601}},
{{9'sd202, 12'sd-1762, 12'sd1497}, {12'sd-1490, 11'sd711, 13'sd2871}, {10'sd-334, 12'sd1566, 13'sd2417}},
{{14'sd4687, 13'sd2182, 14'sd-7742}, {13'sd3683, 12'sd-1141, 14'sd-4225}, {12'sd-1102, 12'sd1729, 11'sd-613}},
{{8'sd-105, 10'sd-459, 8'sd125}, {12'sd2018, 13'sd2486, 10'sd-492}, {13'sd2320, 12'sd-1191, 12'sd-1157}},
{{13'sd-2182, 11'sd761, 13'sd2380}, {13'sd2711, 11'sd515, 11'sd553}, {11'sd-886, 11'sd-819, 12'sd1228}},
{{13'sd3243, 13'sd3509, 13'sd3580}, {12'sd-1442, 11'sd800, 11'sd675}, {13'sd-2447, 13'sd-2594, 13'sd-2322}},
{{13'sd2386, 13'sd2505, 13'sd-2284}, {7'sd-36, 12'sd1029, 6'sd28}, {13'sd2139, 10'sd276, 13'sd-2496}},
{{13'sd-2978, 11'sd658, 7'sd-40}, {11'sd-796, 12'sd1874, 13'sd2471}, {12'sd1506, 8'sd-77, 13'sd-2372}},
{{7'sd43, 11'sd1012, 12'sd-1857}, {12'sd1460, 13'sd-2055, 12'sd1062}, {7'sd-62, 8'sd-115, 13'sd2178}},
{{11'sd784, 10'sd360, 12'sd-1958}, {13'sd2588, 13'sd-2067, 12'sd-1360}, {12'sd1835, 5'sd-8, 10'sd403}},
{{9'sd217, 12'sd-1217, 13'sd-2780}, {12'sd1894, 13'sd2098, 6'sd-23}, {13'sd2328, 12'sd1757, 13'sd-2177}},
{{12'sd1825, 13'sd-2323, 11'sd927}, {11'sd627, 12'sd-1598, 12'sd-1213}, {12'sd-1959, 11'sd-539, 12'sd-1724}},
{{11'sd947, 12'sd-1665, 11'sd-603}, {12'sd-2013, 12'sd-1827, 13'sd2073}, {13'sd-2464, 12'sd1025, 12'sd-1191}},
{{13'sd2325, 10'sd422, 12'sd1164}, {13'sd-2165, 13'sd2236, 8'sd125}, {6'sd-20, 12'sd-1725, 12'sd-1304}},
{{13'sd-3827, 13'sd-2361, 8'sd64}, {14'sd-4549, 11'sd-644, 12'sd1215}, {14'sd-4282, 9'sd-135, 12'sd1169}},
{{11'sd-753, 12'sd1515, 13'sd-3373}, {11'sd784, 12'sd1094, 11'sd896}, {13'sd-2078, 13'sd-2279, 13'sd-3093}},
{{12'sd-1557, 13'sd2550, 13'sd-3193}, {12'sd-1772, 12'sd-1414, 11'sd702}, {12'sd-1527, 12'sd-1637, 10'sd283}},
{{13'sd-2504, 12'sd-1514, 13'sd2669}, {12'sd-1190, 12'sd1686, 11'sd-582}, {12'sd1740, 11'sd781, 11'sd896}},
{{12'sd-1943, 13'sd2155, 8'sd-80}, {12'sd1455, 12'sd-2039, 12'sd1552}, {7'sd-35, 9'sd-183, 12'sd-1089}},
{{13'sd2058, 13'sd2089, 13'sd-2592}, {11'sd-691, 13'sd2831, 12'sd-1672}, {11'sd-922, 11'sd-1011, 12'sd1094}},
{{10'sd463, 9'sd-239, 12'sd1387}, {12'sd-1582, 13'sd2715, 12'sd1068}, {11'sd-566, 11'sd-632, 12'sd-1451}},
{{13'sd3665, 12'sd1417, 11'sd-854}, {11'sd-868, 13'sd2666, 10'sd-429}, {12'sd1076, 13'sd-2395, 13'sd-2500}},
{{13'sd2386, 13'sd2357, 9'sd186}, {13'sd3659, 12'sd1327, 11'sd686}, {13'sd3549, 11'sd778, 11'sd-733}},
{{12'sd1563, 13'sd-2219, 13'sd-2453}, {13'sd-2385, 7'sd-39, 13'sd2173}, {11'sd800, 13'sd-2223, 12'sd1379}},
{{12'sd-1360, 13'sd-3605, 13'sd-2157}, {13'sd-4040, 12'sd-1110, 13'sd-3851}, {13'sd-2674, 13'sd2855, 7'sd32}},
{{12'sd-1177, 12'sd-1483, 12'sd-1049}, {13'sd-2354, 11'sd-728, 13'sd2469}, {13'sd2159, 11'sd585, 11'sd-788}},
{{12'sd-1187, 13'sd2058, 13'sd2245}, {10'sd448, 9'sd178, 11'sd517}, {13'sd2119, 10'sd-278, 12'sd-1249}},
{{13'sd2122, 8'sd-105, 12'sd1876}, {10'sd-474, 12'sd-1065, 12'sd-1193}, {12'sd1875, 13'sd2448, 12'sd-1272}},
{{13'sd2595, 12'sd1075, 13'sd3930}, {12'sd1658, 12'sd-1583, 6'sd17}, {12'sd-1913, 11'sd890, 12'sd1435}},
{{13'sd2248, 13'sd2567, 11'sd728}, {10'sd282, 12'sd-1827, 12'sd1276}, {13'sd-2827, 12'sd1867, 11'sd-906}},
{{12'sd-1849, 10'sd470, 11'sd762}, {13'sd-2874, 12'sd-2046, 13'sd-2746}, {13'sd-2350, 11'sd-995, 12'sd1657}},
{{11'sd901, 9'sd141, 12'sd1349}, {11'sd941, 11'sd963, 14'sd5202}, {12'sd1830, 9'sd204, 14'sd5167}},
{{13'sd-2374, 12'sd1126, 12'sd-1350}, {13'sd-3006, 13'sd2067, 13'sd-2861}, {12'sd-1261, 13'sd2290, 12'sd1813}},
{{13'sd-2100, 11'sd-724, 11'sd-913}, {10'sd354, 11'sd-1020, 12'sd-1252}, {13'sd2195, 12'sd2045, 5'sd-13}},
{{12'sd1203, 13'sd-3335, 12'sd-1088}, {12'sd-1081, 12'sd1343, 12'sd-1146}, {13'sd-2993, 12'sd1463, 13'sd-2095}},
{{13'sd2973, 11'sd1010, 12'sd1648}, {13'sd2570, 11'sd972, 12'sd-1184}, {12'sd1891, 12'sd-1364, 12'sd-1569}},
{{9'sd-255, 12'sd1469, 11'sd-830}, {11'sd-702, 9'sd219, 12'sd1677}, {13'sd-2335, 10'sd-461, 12'sd1829}},
{{11'sd-883, 11'sd518, 11'sd-899}, {10'sd507, 12'sd-1214, 13'sd-2052}, {13'sd2727, 12'sd1521, 12'sd1863}},
{{13'sd3010, 13'sd3461, 12'sd1229}, {13'sd2362, 12'sd1562, 11'sd-618}, {11'sd-562, 13'sd2158, 9'sd-232}},
{{11'sd837, 12'sd-1862, 13'sd2354}, {12'sd-1060, 13'sd-2541, 12'sd-1498}, {11'sd812, 12'sd-1871, 12'sd1159}},
{{12'sd-1097, 12'sd-1812, 13'sd-3833}, {6'sd-24, 9'sd188, 11'sd1012}, {11'sd559, 12'sd1193, 8'sd77}},
{{12'sd-1285, 10'sd381, 10'sd-328}, {13'sd2132, 11'sd-794, 13'sd2763}, {12'sd1720, 11'sd722, 13'sd2510}},
{{12'sd-1040, 12'sd1888, 12'sd-1867}, {11'sd675, 10'sd-310, 11'sd-671}, {13'sd-3956, 9'sd180, 12'sd-1517}},
{{11'sd-827, 13'sd-2311, 12'sd1266}, {13'sd-3091, 11'sd-948, 13'sd3036}, {13'sd2592, 12'sd-1374, 12'sd-1200}},
{{12'sd-1521, 11'sd786, 12'sd2044}, {13'sd2414, 12'sd1699, 10'sd494}, {10'sd-488, 13'sd-3360, 11'sd-1022}},
{{10'sd495, 11'sd-808, 12'sd1575}, {12'sd-1414, 12'sd1917, 11'sd-732}, {12'sd-1834, 11'sd676, 13'sd-2416}},
{{11'sd-722, 11'sd675, 12'sd1759}, {12'sd-1379, 13'sd-2125, 12'sd1908}, {13'sd2208, 10'sd-316, 12'sd1992}},
{{13'sd3523, 13'sd2633, 9'sd128}, {9'sd-181, 13'sd2089, 13'sd-4093}, {13'sd-2102, 10'sd-394, 14'sd-5072}},
{{8'sd-125, 13'sd2394, 12'sd1966}, {11'sd860, 12'sd-1344, 13'sd2327}, {10'sd294, 10'sd-434, 11'sd944}},
{{11'sd-524, 12'sd-1605, 13'sd-2545}, {11'sd-546, 10'sd499, 11'sd848}, {8'sd74, 12'sd-1420, 13'sd-2097}},
{{12'sd1330, 12'sd1983, 13'sd3883}, {11'sd554, 10'sd-441, 13'sd3074}, {11'sd-659, 12'sd1579, 8'sd81}},
{{12'sd-2029, 10'sd393, 13'sd-2900}, {11'sd514, 12'sd-1396, 13'sd-2606}, {6'sd-22, 11'sd-721, 10'sd298}}},
{
{{13'sd-2593, 11'sd667, 12'sd-1861}, {12'sd1235, 13'sd2412, 12'sd2035}, {11'sd-816, 12'sd-1749, 12'sd1273}},
{{11'sd644, 10'sd471, 11'sd-758}, {12'sd1336, 11'sd991, 9'sd-214}, {13'sd2239, 12'sd-1555, 13'sd2439}},
{{13'sd2567, 13'sd-2366, 10'sd-358}, {12'sd-1823, 13'sd2075, 11'sd992}, {12'sd-1333, 13'sd-2527, 10'sd-496}},
{{13'sd-2312, 11'sd910, 11'sd966}, {13'sd2342, 10'sd389, 13'sd-2646}, {12'sd1245, 12'sd-1680, 12'sd-1643}},
{{12'sd-1319, 13'sd-2481, 13'sd-2537}, {12'sd-1330, 13'sd2187, 13'sd2573}, {11'sd685, 10'sd-474, 12'sd-1583}},
{{7'sd-45, 12'sd-1879, 13'sd3085}, {11'sd545, 12'sd-1601, 13'sd3022}, {11'sd-935, 12'sd-1616, 11'sd727}},
{{13'sd2125, 11'sd986, 12'sd1544}, {12'sd1413, 12'sd-1306, 12'sd-1395}, {13'sd-2157, 6'sd-26, 11'sd901}},
{{12'sd1338, 8'sd-108, 11'sd-950}, {12'sd-1944, 13'sd2230, 9'sd-241}, {12'sd-1515, 13'sd-2555, 11'sd-862}},
{{13'sd-2556, 7'sd41, 7'sd58}, {12'sd1540, 12'sd-1927, 12'sd1935}, {12'sd-1569, 12'sd1544, 12'sd1494}},
{{12'sd-1718, 9'sd236, 11'sd-625}, {12'sd1706, 12'sd-1163, 12'sd1681}, {10'sd-479, 12'sd-1149, 11'sd-687}},
{{10'sd372, 12'sd1219, 13'sd-2328}, {12'sd1163, 10'sd-293, 12'sd-1224}, {11'sd-896, 12'sd1537, 12'sd-1759}},
{{11'sd-549, 13'sd-2392, 12'sd-1520}, {10'sd-338, 8'sd-126, 10'sd314}, {13'sd2063, 12'sd-1773, 10'sd403}},
{{13'sd-2235, 13'sd-2598, 13'sd-2240}, {12'sd-1469, 12'sd1372, 13'sd-2667}, {13'sd2582, 12'sd1385, 11'sd740}},
{{12'sd-1403, 12'sd-1288, 12'sd-1882}, {13'sd-2519, 13'sd-2211, 11'sd944}, {12'sd2016, 11'sd882, 12'sd-1075}},
{{9'sd-192, 6'sd-28, 12'sd-1800}, {13'sd-2465, 13'sd3413, 11'sd678}, {11'sd-872, 9'sd-214, 12'sd-1189}},
{{11'sd-718, 10'sd-363, 12'sd1924}, {12'sd1246, 12'sd-1222, 13'sd-2711}, {9'sd190, 13'sd2309, 12'sd-1278}},
{{11'sd-873, 10'sd369, 12'sd-1593}, {13'sd-2622, 13'sd2083, 13'sd2267}, {13'sd-2160, 13'sd-2240, 11'sd561}},
{{12'sd1585, 12'sd1419, 11'sd-878}, {12'sd1655, 13'sd-2302, 11'sd-639}, {12'sd1880, 12'sd1664, 11'sd813}},
{{12'sd1115, 10'sd-271, 12'sd1568}, {10'sd-467, 10'sd-301, 11'sd850}, {13'sd-2431, 12'sd-1633, 10'sd-400}},
{{12'sd-1783, 12'sd-1228, 12'sd-1373}, {12'sd1451, 12'sd2006, 9'sd247}, {12'sd-1332, 11'sd-1002, 11'sd-1011}},
{{11'sd588, 12'sd-1222, 12'sd-1516}, {13'sd-2931, 12'sd1274, 10'sd462}, {13'sd-2350, 11'sd600, 13'sd-2268}},
{{12'sd1140, 9'sd-140, 12'sd1650}, {12'sd2029, 12'sd-1838, 12'sd1854}, {12'sd-1619, 12'sd-1632, 12'sd-1650}},
{{12'sd1488, 11'sd772, 12'sd1867}, {12'sd1136, 13'sd2690, 13'sd2712}, {11'sd585, 13'sd2422, 12'sd1450}},
{{10'sd-477, 11'sd970, 12'sd-1185}, {10'sd-457, 9'sd-214, 12'sd1734}, {8'sd-124, 13'sd-2411, 12'sd-1926}},
{{12'sd-1351, 13'sd-2221, 10'sd300}, {11'sd-556, 10'sd-391, 11'sd968}, {12'sd-1711, 11'sd582, 13'sd2365}},
{{11'sd-585, 11'sd792, 12'sd1299}, {13'sd2484, 13'sd2765, 11'sd-564}, {12'sd1813, 11'sd-952, 12'sd-1613}},
{{12'sd-1560, 8'sd81, 12'sd1394}, {13'sd-3010, 13'sd-2631, 10'sd315}, {13'sd-3050, 13'sd-3551, 10'sd-409}},
{{13'sd-2442, 9'sd-145, 12'sd-1649}, {13'sd-2128, 13'sd-2397, 11'sd-718}, {10'sd-257, 12'sd-1142, 13'sd-2137}},
{{13'sd2275, 11'sd-1020, 13'sd-2179}, {12'sd-1763, 11'sd538, 12'sd1698}, {12'sd-1247, 11'sd634, 11'sd-651}},
{{13'sd-2942, 12'sd-1401, 10'sd344}, {11'sd814, 12'sd-1956, 12'sd1385}, {13'sd2322, 12'sd1558, 11'sd-686}},
{{12'sd-1157, 12'sd1059, 11'sd-721}, {13'sd-2156, 10'sd-301, 8'sd100}, {12'sd1371, 13'sd2473, 12'sd1119}},
{{11'sd-919, 13'sd-2243, 13'sd2681}, {11'sd-755, 12'sd-1571, 12'sd-1159}, {12'sd2032, 10'sd-389, 11'sd590}},
{{6'sd16, 11'sd-554, 11'sd-573}, {12'sd-1887, 6'sd26, 11'sd843}, {10'sd-350, 13'sd2142, 7'sd38}},
{{13'sd2587, 13'sd-2477, 13'sd-2088}, {12'sd1670, 13'sd2365, 11'sd529}, {12'sd-2004, 12'sd-1370, 11'sd-721}},
{{13'sd-2853, 13'sd2234, 11'sd-1014}, {12'sd-2046, 12'sd1175, 13'sd-2518}, {13'sd-2676, 12'sd1900, 13'sd-2551}},
{{11'sd915, 12'sd-1610, 7'sd-40}, {11'sd633, 10'sd-413, 12'sd1237}, {9'sd243, 13'sd-2342, 10'sd474}},
{{9'sd-167, 11'sd-549, 12'sd1841}, {12'sd-1601, 7'sd-57, 13'sd-2050}, {7'sd-48, 12'sd-1609, 12'sd-1834}},
{{10'sd302, 11'sd568, 13'sd-2196}, {11'sd707, 13'sd-2651, 11'sd-708}, {12'sd-1339, 12'sd1700, 11'sd-918}},
{{12'sd-1197, 12'sd-1397, 12'sd1385}, {11'sd920, 13'sd-2665, 12'sd-1646}, {12'sd1625, 10'sd412, 9'sd-205}},
{{12'sd1436, 10'sd-342, 10'sd-443}, {12'sd-1541, 13'sd2202, 13'sd2187}, {12'sd1932, 9'sd131, 9'sd213}},
{{12'sd1795, 11'sd723, 9'sd228}, {12'sd-1661, 13'sd-2480, 11'sd553}, {12'sd-1853, 11'sd-755, 10'sd-477}},
{{11'sd-716, 13'sd2277, 10'sd371}, {11'sd-770, 12'sd-1737, 11'sd753}, {9'sd220, 10'sd390, 11'sd-548}},
{{13'sd-2171, 10'sd-470, 9'sd-131}, {13'sd2502, 12'sd-1355, 12'sd-1586}, {13'sd-2149, 12'sd-1127, 13'sd-2056}},
{{11'sd949, 13'sd-3081, 13'sd-2782}, {13'sd3320, 11'sd-733, 13'sd-2338}, {11'sd-845, 13'sd-2920, 10'sd325}},
{{11'sd695, 13'sd2470, 12'sd1194}, {12'sd-1296, 13'sd2121, 9'sd-235}, {8'sd-64, 10'sd-371, 7'sd63}},
{{13'sd2321, 13'sd2667, 12'sd1360}, {13'sd2365, 12'sd-1587, 13'sd2129}, {11'sd-809, 12'sd-1597, 10'sd387}},
{{12'sd1222, 13'sd2122, 11'sd762}, {12'sd-1178, 12'sd-1268, 13'sd-2343}, {11'sd565, 11'sd-515, 13'sd-2323}},
{{13'sd-3053, 10'sd434, 9'sd-211}, {8'sd-120, 12'sd-1742, 12'sd1460}, {12'sd1545, 12'sd-1688, 12'sd2013}},
{{12'sd-1414, 9'sd222, 12'sd1612}, {11'sd822, 9'sd-190, 13'sd-2185}, {12'sd-1210, 13'sd2153, 12'sd1249}},
{{12'sd-1197, 13'sd2659, 10'sd422}, {12'sd-1116, 13'sd-2055, 7'sd49}, {12'sd1703, 13'sd2716, 9'sd148}},
{{11'sd571, 12'sd1544, 9'sd223}, {12'sd1413, 12'sd1362, 8'sd86}, {12'sd1372, 12'sd2004, 8'sd-115}},
{{11'sd701, 12'sd-1582, 5'sd8}, {11'sd-702, 11'sd-643, 13'sd2554}, {12'sd-1287, 13'sd-2517, 11'sd685}},
{{11'sd779, 13'sd2246, 12'sd-1660}, {12'sd-1954, 13'sd3497, 10'sd510}, {13'sd-2236, 12'sd1658, 12'sd-1307}},
{{12'sd-1263, 13'sd2487, 12'sd-1474}, {11'sd833, 10'sd263, 13'sd-2553}, {11'sd659, 11'sd676, 12'sd-1815}},
{{11'sd646, 12'sd1657, 13'sd-3128}, {12'sd1859, 11'sd-692, 12'sd1514}, {13'sd-2770, 12'sd1875, 13'sd2107}},
{{13'sd-2081, 12'sd1864, 12'sd-1416}, {13'sd2249, 12'sd-1890, 12'sd1866}, {9'sd-173, 12'sd1466, 13'sd2412}},
{{10'sd-398, 12'sd-1246, 12'sd-2012}, {12'sd1628, 12'sd-1428, 10'sd318}, {12'sd-2032, 11'sd-687, 12'sd-1962}},
{{11'sd1012, 12'sd-2034, 11'sd772}, {12'sd1409, 12'sd-1689, 12'sd1379}, {13'sd-2203, 12'sd1091, 12'sd1026}},
{{13'sd2137, 12'sd-1764, 13'sd-2074}, {12'sd1603, 12'sd-1524, 12'sd1796}, {9'sd245, 12'sd-1578, 11'sd962}},
{{10'sd-276, 12'sd-1311, 13'sd2147}, {12'sd-1889, 12'sd1517, 13'sd2716}, {10'sd-475, 12'sd1168, 10'sd491}},
{{12'sd-1495, 12'sd-1807, 9'sd207}, {12'sd-1918, 11'sd837, 13'sd-2769}, {12'sd1430, 13'sd2604, 11'sd598}},
{{12'sd1802, 9'sd248, 13'sd-2181}, {12'sd-1467, 11'sd-514, 13'sd-2086}, {13'sd2060, 12'sd1340, 11'sd-801}},
{{9'sd-132, 10'sd481, 9'sd-130}, {12'sd1415, 12'sd-1492, 12'sd1427}, {13'sd-2501, 12'sd1994, 10'sd-293}},
{{12'sd-1789, 9'sd-176, 12'sd-1943}, {13'sd2876, 12'sd1420, 11'sd977}, {12'sd1686, 13'sd2209, 11'sd-600}}},
{
{{12'sd-1927, 12'sd-1321, 13'sd-2173}, {11'sd886, 11'sd547, 12'sd-1828}, {12'sd1601, 10'sd511, 12'sd-1208}},
{{12'sd1244, 12'sd-1320, 13'sd2427}, {11'sd-576, 12'sd1045, 13'sd-2663}, {7'sd37, 13'sd-2610, 12'sd-1858}},
{{11'sd-872, 12'sd1419, 10'sd-335}, {10'sd438, 12'sd-1448, 13'sd-2495}, {12'sd-1742, 8'sd71, 12'sd1608}},
{{9'sd175, 13'sd2586, 12'sd-1961}, {11'sd732, 11'sd561, 12'sd-1781}, {11'sd-649, 12'sd1433, 9'sd151}},
{{11'sd538, 11'sd-701, 12'sd-1724}, {13'sd3870, 11'sd1017, 11'sd-843}, {8'sd82, 13'sd3045, 13'sd3286}},
{{13'sd-2470, 11'sd-696, 13'sd-2401}, {13'sd-2170, 12'sd-1895, 12'sd-1330}, {13'sd2373, 12'sd1919, 12'sd-1291}},
{{13'sd2059, 6'sd-24, 13'sd2862}, {13'sd2426, 12'sd-1998, 13'sd2204}, {13'sd2761, 12'sd-1636, 13'sd2614}},
{{12'sd1892, 12'sd1615, 11'sd727}, {13'sd2532, 10'sd-306, 12'sd-1664}, {10'sd-446, 13'sd2353, 13'sd-2346}},
{{12'sd-1338, 13'sd2510, 13'sd2414}, {11'sd-546, 13'sd-2663, 11'sd627}, {11'sd793, 12'sd1041, 7'sd-55}},
{{12'sd1249, 10'sd-477, 12'sd-1958}, {12'sd-1555, 13'sd3437, 10'sd-442}, {12'sd-1643, 13'sd2974, 9'sd154}},
{{11'sd-739, 11'sd695, 13'sd2509}, {13'sd-2253, 13'sd2682, 12'sd1828}, {11'sd981, 9'sd144, 12'sd-1520}},
{{9'sd202, 12'sd1423, 11'sd904}, {12'sd1182, 13'sd2238, 9'sd-187}, {12'sd1419, 11'sd-558, 10'sd491}},
{{12'sd1938, 12'sd-1836, 13'sd-2264}, {10'sd-428, 13'sd2808, 12'sd-1812}, {12'sd-1987, 10'sd335, 13'sd2753}},
{{11'sd-998, 13'sd2570, 11'sd-943}, {12'sd-1546, 7'sd60, 11'sd649}, {13'sd-2135, 10'sd287, 13'sd-2168}},
{{13'sd-3243, 12'sd-1186, 11'sd-769}, {12'sd-1507, 12'sd-1401, 12'sd1822}, {12'sd-1789, 11'sd965, 11'sd592}},
{{11'sd599, 11'sd612, 10'sd507}, {12'sd1043, 9'sd-185, 12'sd-1058}, {12'sd-1735, 12'sd1560, 12'sd1663}},
{{9'sd-239, 11'sd831, 11'sd826}, {11'sd977, 10'sd486, 9'sd-239}, {12'sd-1065, 12'sd-1105, 11'sd976}},
{{12'sd-1738, 12'sd-1046, 12'sd-1783}, {13'sd2185, 12'sd-1552, 12'sd1246}, {10'sd355, 12'sd-1285, 12'sd1771}},
{{12'sd1699, 9'sd225, 11'sd945}, {12'sd-1090, 10'sd273, 12'sd1093}, {13'sd-2313, 12'sd1811, 13'sd2235}},
{{12'sd1773, 13'sd-2240, 13'sd2519}, {12'sd1668, 12'sd-1045, 6'sd17}, {12'sd-1383, 12'sd-1467, 12'sd-1469}},
{{12'sd-1431, 10'sd460, 12'sd-1927}, {12'sd1481, 12'sd-1292, 12'sd1374}, {10'sd-448, 13'sd-2600, 11'sd-529}},
{{11'sd595, 13'sd-2539, 8'sd-81}, {13'sd2202, 13'sd2519, 12'sd1334}, {11'sd733, 11'sd564, 12'sd-1070}},
{{13'sd2529, 11'sd979, 8'sd-109}, {13'sd3056, 13'sd3067, 12'sd-1350}, {12'sd-1537, 9'sd140, 13'sd-2156}},
{{12'sd-1796, 12'sd1383, 12'sd-1108}, {10'sd-430, 13'sd-2228, 12'sd-1573}, {12'sd-1861, 13'sd2188, 8'sd73}},
{{13'sd2619, 12'sd-1729, 12'sd1833}, {12'sd-1322, 13'sd-2243, 9'sd233}, {13'sd-2496, 11'sd-616, 12'sd1732}},
{{9'sd-252, 13'sd2203, 12'sd-1611}, {12'sd-1602, 12'sd-1266, 13'sd-2578}, {13'sd2258, 12'sd1266, 9'sd-212}},
{{12'sd-1206, 13'sd-2184, 11'sd908}, {12'sd1574, 10'sd496, 13'sd-3191}, {12'sd-1649, 12'sd-1461, 13'sd-3263}},
{{12'sd-1348, 11'sd642, 12'sd-1825}, {13'sd2529, 10'sd420, 12'sd-2010}, {11'sd-1014, 12'sd1628, 12'sd-1609}},
{{12'sd1871, 7'sd-53, 11'sd745}, {9'sd-160, 12'sd1205, 9'sd-203}, {12'sd1736, 12'sd1212, 12'sd1359}},
{{8'sd85, 13'sd-2340, 12'sd1178}, {13'sd-2392, 12'sd1993, 12'sd1431}, {13'sd-2624, 10'sd-335, 11'sd-971}},
{{11'sd-773, 13'sd-2180, 12'sd1642}, {12'sd-1866, 13'sd-2196, 12'sd1161}, {12'sd1569, 13'sd-2161, 12'sd-1024}},
{{13'sd2223, 10'sd-391, 12'sd-1671}, {12'sd1838, 13'sd-2608, 11'sd-745}, {13'sd2650, 12'sd-1402, 12'sd-1642}},
{{13'sd2797, 13'sd-2882, 13'sd-2577}, {10'sd-439, 11'sd-862, 11'sd-889}, {12'sd-1315, 10'sd-299, 13'sd2064}},
{{11'sd-707, 9'sd209, 10'sd388}, {12'sd-1180, 9'sd163, 11'sd887}, {12'sd1523, 13'sd-2803, 11'sd862}},
{{12'sd-1992, 13'sd-3145, 12'sd-1278}, {13'sd-2445, 10'sd456, 13'sd-2191}, {11'sd767, 13'sd-3141, 12'sd1448}},
{{11'sd-806, 13'sd-2300, 11'sd-904}, {13'sd-2224, 10'sd-497, 12'sd1581}, {12'sd-1219, 13'sd2654, 12'sd2042}},
{{11'sd750, 14'sd-4782, 11'sd-568}, {1'sd0, 9'sd-146, 8'sd84}, {13'sd-2914, 14'sd-4423, 13'sd-2938}},
{{13'sd2684, 12'sd-1690, 12'sd-1780}, {12'sd1179, 12'sd1900, 12'sd1693}, {13'sd3072, 13'sd2153, 9'sd-222}},
{{10'sd360, 12'sd-1570, 12'sd1965}, {11'sd-895, 12'sd-1766, 8'sd-110}, {11'sd-528, 12'sd-1084, 13'sd-2378}},
{{9'sd239, 12'sd-1106, 5'sd-9}, {13'sd2384, 13'sd-2108, 9'sd210}, {11'sd779, 12'sd-1406, 12'sd1860}},
{{12'sd1409, 13'sd2238, 11'sd683}, {13'sd-2162, 12'sd1466, 12'sd-1681}, {11'sd-634, 11'sd877, 12'sd-2047}},
{{12'sd-1598, 11'sd-970, 8'sd-84}, {9'sd236, 13'sd3363, 13'sd-2109}, {12'sd1637, 13'sd2790, 12'sd1026}},
{{11'sd532, 12'sd1050, 13'sd2474}, {8'sd-99, 12'sd1937, 12'sd-1484}, {10'sd-359, 10'sd-484, 12'sd1189}},
{{12'sd-1207, 13'sd2583, 13'sd-3352}, {12'sd1048, 13'sd-2548, 13'sd2160}, {12'sd-1310, 11'sd1008, 10'sd-313}},
{{12'sd-1296, 12'sd1184, 12'sd-1952}, {12'sd1177, 12'sd1657, 12'sd-1707}, {13'sd-2332, 13'sd-2590, 13'sd-2540}},
{{8'sd-125, 12'sd-1292, 12'sd-1934}, {12'sd1148, 11'sd980, 11'sd-769}, {13'sd2308, 13'sd-2461, 13'sd2302}},
{{13'sd-3032, 12'sd-1423, 13'sd2143}, {11'sd-579, 13'sd-3316, 11'sd794}, {12'sd-1950, 13'sd-2782, 10'sd298}},
{{9'sd163, 13'sd2308, 11'sd-869}, {12'sd1995, 13'sd2064, 12'sd-1535}, {12'sd1125, 10'sd-491, 10'sd401}},
{{12'sd1394, 11'sd733, 13'sd2058}, {13'sd-3215, 12'sd-1676, 13'sd-2393}, {13'sd-2318, 13'sd-3202, 13'sd-2911}},
{{13'sd2700, 13'sd-3038, 11'sd-879}, {10'sd292, 11'sd-903, 12'sd1128}, {10'sd-329, 11'sd-657, 12'sd-1888}},
{{5'sd-10, 11'sd837, 11'sd630}, {13'sd2315, 13'sd2782, 13'sd2696}, {13'sd-2351, 11'sd854, 11'sd-734}},
{{11'sd1000, 13'sd2079, 8'sd121}, {9'sd-167, 13'sd2637, 12'sd-1509}, {13'sd2825, 12'sd-1254, 12'sd1186}},
{{7'sd35, 13'sd2736, 10'sd354}, {8'sd-110, 11'sd-751, 12'sd1299}, {11'sd-708, 13'sd2302, 10'sd-375}},
{{11'sd-677, 10'sd286, 7'sd-61}, {7'sd50, 12'sd1680, 11'sd-875}, {11'sd-665, 13'sd-2080, 11'sd834}},
{{13'sd2310, 13'sd-2108, 13'sd2847}, {10'sd321, 12'sd-1781, 12'sd-1929}, {12'sd-1171, 11'sd-931, 13'sd2495}},
{{11'sd871, 13'sd-3267, 13'sd2335}, {10'sd307, 13'sd-3077, 11'sd717}, {11'sd-824, 10'sd-507, 12'sd-1999}},
{{12'sd1164, 13'sd3037, 11'sd-912}, {13'sd2095, 12'sd1783, 12'sd-1829}, {14'sd4544, 10'sd509, 13'sd2672}},
{{4'sd-6, 13'sd-2421, 12'sd-1131}, {12'sd1296, 12'sd-1414, 12'sd-1740}, {12'sd-1627, 9'sd-166, 12'sd1940}},
{{11'sd738, 12'sd1350, 11'sd1003}, {12'sd1772, 12'sd-1701, 11'sd-547}, {13'sd2108, 11'sd950, 12'sd1942}},
{{13'sd-3149, 13'sd-2185, 12'sd1551}, {11'sd875, 12'sd1109, 13'sd2553}, {12'sd-1344, 7'sd-49, 10'sd378}},
{{13'sd2401, 10'sd460, 12'sd1730}, {12'sd-1536, 12'sd1863, 12'sd-1102}, {13'sd2156, 12'sd-1388, 12'sd-1939}},
{{12'sd-1480, 13'sd-2271, 12'sd1824}, {13'sd2150, 10'sd-443, 13'sd-2769}, {12'sd1159, 12'sd1174, 12'sd-1282}},
{{13'sd-2140, 11'sd-849, 12'sd1244}, {12'sd-1359, 10'sd373, 10'sd-476}, {7'sd45, 11'sd-998, 11'sd650}},
{{12'sd1445, 11'sd-842, 11'sd-543}, {13'sd-2719, 10'sd313, 12'sd1511}, {11'sd638, 12'sd1761, 12'sd1061}}},
{
{{12'sd1722, 11'sd-611, 11'sd-918}, {12'sd1879, 13'sd-2355, 10'sd-459}, {7'sd57, 9'sd-201, 13'sd3006}},
{{13'sd-2463, 13'sd2090, 11'sd-817}, {13'sd2278, 12'sd1651, 10'sd374}, {11'sd-914, 9'sd-215, 11'sd-772}},
{{10'sd313, 12'sd1094, 10'sd270}, {11'sd-798, 12'sd-1707, 13'sd2692}, {13'sd-2685, 12'sd1389, 12'sd-1227}},
{{11'sd567, 12'sd-1579, 12'sd-1437}, {12'sd-1395, 12'sd-1267, 13'sd2162}, {12'sd1737, 12'sd-1570, 12'sd-1602}},
{{12'sd-1514, 12'sd-1546, 13'sd3505}, {13'sd2795, 13'sd3154, 14'sd4591}, {10'sd304, 12'sd1784, 13'sd2801}},
{{12'sd-1597, 13'sd2761, 10'sd412}, {12'sd1193, 13'sd3210, 13'sd3176}, {11'sd578, 13'sd3689, 13'sd2056}},
{{12'sd1834, 13'sd2903, 13'sd3369}, {13'sd-2540, 13'sd2221, 11'sd-546}, {12'sd-1692, 11'sd516, 11'sd530}},
{{10'sd-485, 9'sd-248, 13'sd2270}, {10'sd400, 11'sd-568, 11'sd784}, {12'sd-1604, 12'sd1311, 13'sd-2090}},
{{11'sd-983, 13'sd-2309, 11'sd909}, {12'sd-1097, 12'sd-1409, 13'sd-2124}, {12'sd-1625, 11'sd724, 13'sd-2273}},
{{11'sd-592, 10'sd469, 11'sd-513}, {5'sd-13, 12'sd-1198, 10'sd280}, {12'sd-2035, 10'sd445, 13'sd2626}},
{{13'sd-3147, 8'sd75, 12'sd-1902}, {10'sd317, 11'sd-872, 12'sd1142}, {13'sd-2507, 12'sd-1931, 12'sd-1063}},
{{12'sd-1033, 12'sd-1320, 12'sd-1262}, {13'sd2668, 12'sd-1770, 13'sd-2553}, {13'sd-2091, 13'sd2444, 9'sd165}},
{{10'sd348, 8'sd-113, 12'sd1706}, {13'sd-2094, 10'sd-266, 12'sd1939}, {12'sd-1556, 12'sd-2000, 12'sd1216}},
{{9'sd205, 13'sd-2096, 13'sd2232}, {11'sd708, 13'sd-2559, 12'sd-1796}, {12'sd-1925, 13'sd-2873, 11'sd-629}},
{{12'sd-1252, 12'sd2008, 11'sd-1004}, {11'sd539, 13'sd-3431, 13'sd-2388}, {12'sd-1375, 11'sd-1005, 12'sd-1405}},
{{12'sd1326, 8'sd-92, 10'sd411}, {11'sd-831, 9'sd186, 12'sd1203}, {12'sd1117, 13'sd2877, 9'sd190}},
{{13'sd2621, 12'sd1678, 13'sd-2660}, {11'sd960, 12'sd-1178, 12'sd1389}, {11'sd875, 12'sd1384, 10'sd511}},
{{12'sd-1268, 9'sd232, 11'sd-592}, {12'sd1052, 12'sd1989, 11'sd857}, {12'sd-1248, 12'sd1742, 11'sd-763}},
{{13'sd-2561, 13'sd2509, 12'sd1313}, {12'sd1492, 11'sd922, 12'sd1265}, {11'sd-631, 11'sd-903, 10'sd257}},
{{13'sd2452, 12'sd1988, 10'sd-364}, {12'sd-1095, 11'sd-711, 13'sd-2240}, {12'sd1309, 13'sd-2433, 12'sd-1595}},
{{10'sd435, 12'sd-1954, 8'sd-102}, {9'sd-198, 12'sd1238, 12'sd-1296}, {12'sd1073, 12'sd-1060, 11'sd-619}},
{{12'sd1111, 12'sd1289, 13'sd-2253}, {11'sd726, 12'sd1392, 11'sd838}, {13'sd2504, 13'sd2195, 13'sd2070}},
{{11'sd-928, 12'sd1434, 12'sd1545}, {13'sd2230, 13'sd2409, 10'sd284}, {11'sd562, 12'sd1828, 13'sd-2148}},
{{7'sd-62, 11'sd743, 11'sd-737}, {10'sd-339, 12'sd-1861, 12'sd-1948}, {11'sd-1012, 10'sd504, 10'sd327}},
{{11'sd-517, 13'sd-2157, 12'sd-2045}, {12'sd-1893, 6'sd-21, 13'sd-2210}, {12'sd1947, 11'sd934, 13'sd-2554}},
{{13'sd-2818, 12'sd-1078, 12'sd-1514}, {13'sd2390, 11'sd-660, 13'sd2888}, {13'sd2172, 13'sd2294, 10'sd-482}},
{{12'sd-1969, 11'sd591, 13'sd2372}, {11'sd978, 13'sd-2481, 8'sd-124}, {12'sd-1681, 11'sd1016, 8'sd72}},
{{13'sd2782, 12'sd1787, 12'sd-1363}, {8'sd-79, 13'sd-2435, 12'sd1790}, {13'sd-2705, 11'sd741, 12'sd1155}},
{{13'sd-2087, 12'sd-1922, 10'sd307}, {13'sd-3250, 13'sd2071, 10'sd421}, {11'sd-801, 11'sd-786, 10'sd-486}},
{{12'sd1282, 11'sd515, 11'sd-603}, {12'sd-1547, 13'sd-2517, 12'sd1526}, {13'sd-2617, 13'sd-2219, 12'sd1522}},
{{12'sd-1645, 12'sd-1289, 11'sd-671}, {11'sd517, 12'sd1246, 13'sd-2382}, {11'sd-923, 13'sd2732, 9'sd-241}},
{{11'sd-617, 12'sd2044, 12'sd1918}, {12'sd1559, 13'sd-2291, 13'sd-2062}, {10'sd299, 13'sd-2225, 13'sd2520}},
{{12'sd-1359, 13'sd2204, 11'sd-801}, {12'sd1815, 12'sd-1385, 12'sd1862}, {11'sd772, 12'sd-1925, 10'sd-420}},
{{10'sd-471, 12'sd-2033, 12'sd1508}, {13'sd-2255, 12'sd-1628, 13'sd-2302}, {12'sd-1538, 13'sd-2910, 11'sd-518}},
{{12'sd2037, 12'sd1767, 12'sd-1853}, {13'sd2385, 6'sd27, 13'sd-2737}, {12'sd1859, 11'sd752, 12'sd-1785}},
{{10'sd-489, 12'sd-1064, 12'sd-1426}, {12'sd1707, 12'sd-1122, 13'sd2065}, {13'sd2554, 13'sd-2634, 12'sd-1323}},
{{13'sd3530, 13'sd2108, 12'sd-1859}, {7'sd-50, 11'sd824, 13'sd-3337}, {12'sd1897, 11'sd-658, 11'sd-813}},
{{13'sd-2071, 8'sd76, 12'sd2017}, {13'sd2117, 12'sd1777, 11'sd-895}, {12'sd1764, 13'sd2645, 11'sd1003}},
{{13'sd-2330, 12'sd1051, 12'sd1588}, {11'sd824, 12'sd2025, 9'sd225}, {13'sd2416, 13'sd-2464, 11'sd568}},
{{7'sd34, 11'sd762, 12'sd1180}, {12'sd1342, 13'sd2586, 13'sd2267}, {12'sd-1889, 12'sd-1332, 13'sd2312}},
{{11'sd-640, 11'sd640, 13'sd2204}, {13'sd2641, 11'sd939, 11'sd-962}, {10'sd-462, 11'sd878, 13'sd2057}},
{{11'sd-616, 11'sd-852, 12'sd1878}, {12'sd1268, 12'sd-1221, 12'sd1692}, {13'sd-2361, 13'sd2592, 12'sd-1303}},
{{11'sd985, 9'sd-241, 11'sd658}, {10'sd-259, 13'sd-2787, 12'sd1548}, {12'sd-1451, 13'sd-2497, 13'sd-3074}},
{{13'sd-2688, 11'sd997, 12'sd-1848}, {12'sd-1848, 13'sd2367, 12'sd-1732}, {12'sd1645, 10'sd-274, 13'sd2912}},
{{11'sd-1006, 13'sd2477, 12'sd-1865}, {13'sd-2815, 12'sd1489, 13'sd2262}, {13'sd2663, 13'sd2099, 12'sd1812}},
{{11'sd813, 12'sd1364, 12'sd-1448}, {13'sd2940, 12'sd-1072, 13'sd-2773}, {12'sd1266, 13'sd2552, 13'sd2555}},
{{11'sd803, 12'sd1843, 12'sd-1928}, {12'sd-1090, 13'sd-2607, 12'sd1263}, {13'sd2458, 11'sd-631, 10'sd-422}},
{{11'sd575, 11'sd-791, 11'sd-782}, {12'sd-1810, 12'sd-1743, 12'sd1492}, {13'sd2914, 13'sd-3329, 13'sd-2778}},
{{12'sd-1506, 10'sd370, 12'sd-1874}, {12'sd1512, 13'sd-2614, 12'sd-1542}, {13'sd2116, 12'sd-1117, 12'sd1120}},
{{13'sd3072, 11'sd-915, 12'sd-1075}, {13'sd3055, 12'sd-2025, 13'sd-2246}, {9'sd174, 11'sd-585, 11'sd986}},
{{12'sd1548, 10'sd-323, 11'sd-925}, {11'sd694, 12'sd1388, 11'sd-839}, {10'sd-455, 11'sd613, 6'sd31}},
{{12'sd1573, 11'sd-944, 10'sd-451}, {10'sd-467, 10'sd-258, 12'sd1794}, {13'sd-2316, 12'sd1412, 12'sd-1744}},
{{12'sd-1144, 13'sd2325, 11'sd-968}, {9'sd-190, 11'sd573, 12'sd-2039}, {5'sd-13, 13'sd-2199, 11'sd807}},
{{10'sd-382, 13'sd2330, 9'sd-232}, {12'sd-1912, 10'sd275, 12'sd-1107}, {13'sd-2252, 12'sd-1147, 11'sd-966}},
{{13'sd3156, 13'sd2959, 13'sd3854}, {12'sd-1076, 12'sd1786, 10'sd406}, {12'sd-1209, 12'sd-1594, 13'sd3793}},
{{11'sd883, 12'sd-1296, 12'sd1812}, {13'sd2825, 10'sd451, 10'sd-259}, {12'sd1456, 12'sd1326, 12'sd-1425}},
{{12'sd1025, 11'sd951, 12'sd1053}, {12'sd-1179, 13'sd2269, 14'sd5619}, {13'sd-2896, 13'sd-3991, 12'sd-1410}},
{{10'sd-344, 11'sd-856, 13'sd-2415}, {5'sd11, 10'sd367, 13'sd2405}, {11'sd-536, 12'sd1595, 11'sd-759}},
{{12'sd1119, 11'sd664, 13'sd2514}, {12'sd-1374, 12'sd1820, 12'sd-1357}, {11'sd569, 13'sd-2726, 13'sd2226}},
{{11'sd679, 7'sd50, 12'sd1290}, {11'sd-684, 12'sd1456, 12'sd-1361}, {12'sd1956, 11'sd868, 11'sd-807}},
{{12'sd-2003, 11'sd-648, 9'sd-186}, {13'sd2431, 12'sd1849, 12'sd-1319}, {10'sd376, 13'sd2788, 12'sd1866}},
{{13'sd2376, 12'sd-1927, 12'sd-1734}, {9'sd-254, 11'sd538, 13'sd2414}, {12'sd1949, 10'sd-432, 12'sd-1042}},
{{13'sd2692, 10'sd441, 10'sd427}, {12'sd-1974, 13'sd2695, 13'sd2487}, {10'sd379, 13'sd3527, 10'sd-374}},
{{12'sd1196, 9'sd221, 13'sd2804}, {13'sd-2664, 11'sd919, 13'sd-2753}, {11'sd-782, 14'sd-4122, 13'sd-2858}}},
{
{{10'sd377, 11'sd752, 11'sd-753}, {8'sd110, 12'sd-1430, 12'sd1249}, {11'sd759, 10'sd-264, 13'sd2508}},
{{11'sd-890, 12'sd1687, 11'sd-914}, {9'sd132, 10'sd379, 13'sd-2375}, {14'sd-4897, 8'sd-106, 12'sd-1328}},
{{3'sd2, 13'sd-3173, 11'sd994}, {11'sd-816, 13'sd2164, 12'sd-1233}, {12'sd1854, 12'sd-1400, 12'sd-1768}},
{{11'sd549, 12'sd1327, 10'sd-349}, {13'sd2989, 11'sd-982, 11'sd630}, {11'sd937, 11'sd676, 12'sd1775}},
{{13'sd-2839, 13'sd-3393, 13'sd-4009}, {10'sd456, 13'sd2258, 11'sd-935}, {10'sd-269, 13'sd2339, 12'sd-1768}},
{{14'sd4720, 13'sd2277, 11'sd700}, {11'sd591, 11'sd935, 14'sd-4687}, {10'sd-436, 12'sd1114, 12'sd1401}},
{{12'sd-1378, 13'sd-3958, 12'sd1403}, {12'sd1782, 11'sd875, 14'sd5271}, {14'sd4293, 14'sd4756, 11'sd624}},
{{12'sd1913, 12'sd-1470, 13'sd-2736}, {12'sd-1940, 13'sd2348, 12'sd1575}, {12'sd-1939, 10'sd-508, 13'sd-2165}},
{{12'sd-1258, 10'sd-444, 11'sd-740}, {12'sd1708, 12'sd-1219, 13'sd2180}, {10'sd262, 12'sd1396, 13'sd-2298}},
{{13'sd-2145, 5'sd10, 13'sd-3721}, {12'sd1286, 12'sd1648, 12'sd-1173}, {12'sd1117, 12'sd-1557, 12'sd-1032}},
{{12'sd-1989, 10'sd-356, 13'sd-2672}, {12'sd1150, 12'sd-1426, 12'sd1786}, {13'sd-3169, 10'sd-313, 13'sd-2664}},
{{13'sd3017, 11'sd-668, 12'sd1580}, {12'sd-1387, 11'sd-988, 9'sd-209}, {9'sd-203, 13'sd-2501, 13'sd-2431}},
{{13'sd-4037, 10'sd358, 12'sd-1951}, {10'sd365, 10'sd-352, 10'sd-447}, {12'sd1949, 11'sd-626, 13'sd2216}},
{{12'sd1384, 7'sd-32, 12'sd-1185}, {13'sd-2978, 12'sd1594, 12'sd-1319}, {12'sd1592, 12'sd-1233, 13'sd-2909}},
{{13'sd3824, 13'sd-2130, 13'sd-2297}, {14'sd6530, 12'sd1045, 13'sd2150}, {15'sd13550, 12'sd1056, 14'sd5590}},
{{14'sd-4242, 11'sd-744, 11'sd-718}, {13'sd-4067, 10'sd480, 13'sd-3080}, {8'sd95, 13'sd-3714, 12'sd1787}},
{{13'sd2130, 11'sd-565, 13'sd-2676}, {10'sd374, 12'sd1948, 10'sd-389}, {13'sd-2260, 13'sd2381, 8'sd88}},
{{12'sd1103, 12'sd-1650, 11'sd-709}, {12'sd2010, 13'sd2154, 12'sd-1385}, {13'sd3145, 11'sd539, 13'sd2611}},
{{13'sd2137, 13'sd2988, 10'sd-297}, {10'sd-396, 11'sd991, 13'sd-2421}, {9'sd-253, 11'sd950, 8'sd81}},
{{12'sd-1214, 12'sd-1160, 13'sd-2565}, {12'sd-1921, 13'sd2332, 13'sd2114}, {4'sd6, 10'sd325, 12'sd1905}},
{{12'sd1454, 9'sd-132, 11'sd-828}, {10'sd381, 13'sd2221, 12'sd-1662}, {13'sd2049, 9'sd-193, 13'sd-2430}},
{{13'sd-2770, 12'sd1538, 12'sd2004}, {9'sd196, 12'sd-1192, 10'sd-360}, {12'sd1038, 12'sd-1585, 12'sd1141}},
{{12'sd-1771, 13'sd-2609, 12'sd1788}, {12'sd-1149, 12'sd-1554, 13'sd-2946}, {8'sd85, 12'sd-1857, 12'sd-1223}},
{{10'sd481, 10'sd331, 12'sd-1085}, {12'sd1060, 11'sd521, 11'sd706}, {13'sd2738, 12'sd1987, 12'sd-1629}},
{{12'sd1250, 10'sd-278, 12'sd1497}, {11'sd-650, 13'sd-2763, 12'sd-1918}, {12'sd-1056, 10'sd384, 12'sd-1185}},
{{12'sd-1487, 12'sd1752, 12'sd1407}, {12'sd-1804, 12'sd-1605, 12'sd-1471}, {12'sd2011, 11'sd876, 13'sd2641}},
{{12'sd1060, 13'sd2188, 12'sd1140}, {13'sd-2957, 11'sd999, 13'sd-2064}, {12'sd-1026, 11'sd547, 13'sd-2413}},
{{12'sd1792, 13'sd-2447, 12'sd1580}, {8'sd-95, 12'sd-1780, 11'sd780}, {14'sd4331, 13'sd3554, 5'sd-9}},
{{13'sd-2123, 13'sd-2629, 12'sd-1161}, {11'sd-721, 13'sd-2432, 6'sd19}, {14'sd-4189, 10'sd296, 11'sd-593}},
{{13'sd3841, 11'sd-830, 13'sd2638}, {13'sd3014, 8'sd86, 13'sd3618}, {13'sd3451, 12'sd1997, 13'sd-2544}},
{{13'sd2708, 12'sd-1826, 9'sd227}, {13'sd-2228, 12'sd-1025, 12'sd-2042}, {11'sd-687, 12'sd-1266, 11'sd709}},
{{12'sd-1691, 12'sd1365, 12'sd-1201}, {12'sd-2032, 12'sd-1828, 11'sd-908}, {14'sd-4105, 13'sd-3097, 11'sd-558}},
{{10'sd-362, 5'sd-13, 9'sd149}, {11'sd952, 11'sd1012, 9'sd-143}, {13'sd2554, 12'sd-1965, 9'sd-167}},
{{11'sd-633, 11'sd-682, 11'sd569}, {13'sd2605, 13'sd2758, 11'sd-740}, {11'sd572, 13'sd2413, 13'sd2175}},
{{11'sd-528, 13'sd-2227, 11'sd-829}, {12'sd-1606, 11'sd-848, 13'sd2835}, {12'sd-1674, 13'sd-2297, 11'sd-754}},
{{12'sd2046, 13'sd-2134, 12'sd-1104}, {8'sd87, 13'sd2181, 12'sd1515}, {11'sd735, 12'sd-1720, 12'sd-1352}},
{{12'sd1802, 13'sd2146, 11'sd516}, {12'sd1687, 13'sd3106, 10'sd-434}, {13'sd2893, 10'sd-307, 12'sd-1200}},
{{11'sd-593, 9'sd234, 12'sd-1567}, {12'sd1889, 12'sd-2019, 12'sd1253}, {12'sd-1436, 13'sd2820, 13'sd3136}},
{{13'sd2504, 10'sd-496, 12'sd1086}, {11'sd-730, 11'sd996, 12'sd-2018}, {12'sd1673, 11'sd-759, 13'sd-2223}},
{{13'sd-2527, 11'sd-782, 12'sd1444}, {11'sd954, 9'sd-131, 11'sd898}, {12'sd-1484, 13'sd-2061, 10'sd488}},
{{12'sd-1078, 10'sd-476, 13'sd-4004}, {13'sd2891, 13'sd2719, 12'sd1654}, {13'sd2997, 9'sd-172, 9'sd-248}},
{{10'sd-404, 12'sd-1731, 12'sd-1594}, {13'sd-3712, 12'sd-1903, 12'sd1154}, {13'sd-3130, 7'sd-44, 10'sd-494}},
{{12'sd1226, 10'sd-323, 14'sd4981}, {13'sd4016, 10'sd-435, 13'sd3412}, {12'sd1484, 12'sd1520, 12'sd-1851}},
{{15'sd-8547, 11'sd-971, 12'sd-1137}, {15'sd-8974, 13'sd-2547, 13'sd-3380}, {15'sd-11480, 14'sd-7013, 14'sd-7609}},
{{12'sd-1267, 6'sd21, 11'sd873}, {13'sd3152, 11'sd-888, 11'sd969}, {12'sd-1360, 12'sd-1142, 12'sd-1406}},
{{13'sd3501, 12'sd-1561, 10'sd-417}, {13'sd-2480, 13'sd2236, 13'sd-2952}, {11'sd916, 13'sd-2088, 13'sd-2058}},
{{8'sd115, 12'sd-1917, 13'sd2288}, {11'sd768, 12'sd1227, 13'sd2674}, {10'sd296, 11'sd928, 12'sd-1414}},
{{12'sd2045, 11'sd553, 13'sd-2171}, {12'sd-1208, 12'sd1172, 13'sd2068}, {13'sd2224, 10'sd-390, 13'sd2136}},
{{14'sd6410, 7'sd-51, 11'sd910}, {13'sd2892, 13'sd3297, 13'sd-2149}, {14'sd5355, 10'sd350, 12'sd-1999}},
{{13'sd2941, 13'sd2406, 9'sd-186}, {13'sd3947, 12'sd1464, 11'sd-550}, {13'sd2911, 13'sd2598, 12'sd-1467}},
{{11'sd897, 12'sd1184, 12'sd-1824}, {11'sd1008, 12'sd-1571, 8'sd-64}, {10'sd417, 12'sd1562, 10'sd277}},
{{12'sd1227, 11'sd935, 11'sd-730}, {12'sd-1131, 13'sd2283, 11'sd860}, {13'sd2349, 13'sd-2386, 12'sd1723}},
{{12'sd1843, 12'sd1146, 10'sd-365}, {10'sd-434, 11'sd839, 8'sd102}, {13'sd3224, 13'sd2694, 12'sd1990}},
{{11'sd773, 12'sd1274, 13'sd2293}, {12'sd-1470, 10'sd-305, 12'sd1435}, {12'sd1347, 12'sd-1659, 13'sd-2681}},
{{13'sd2966, 12'sd1407, 11'sd-565}, {13'sd4082, 12'sd1678, 12'sd-1260}, {14'sd4215, 10'sd449, 13'sd2818}},
{{13'sd2638, 13'sd3024, 13'sd2799}, {11'sd-724, 13'sd2400, 9'sd206}, {12'sd1075, 12'sd-1784, 12'sd-1465}},
{{14'sd-4993, 12'sd-1154, 11'sd-874}, {11'sd-1012, 11'sd-721, 14'sd4669}, {12'sd-1727, 13'sd3247, 10'sd276}},
{{12'sd1778, 9'sd-135, 11'sd-543}, {12'sd1266, 10'sd-495, 12'sd-2046}, {9'sd147, 13'sd-2708, 9'sd-146}},
{{7'sd-38, 13'sd-2232, 12'sd-1053}, {12'sd1169, 6'sd29, 10'sd289}, {10'sd344, 10'sd270, 13'sd2873}},
{{12'sd1483, 13'sd-2663, 12'sd1965}, {13'sd2873, 11'sd-760, 12'sd1326}, {14'sd5713, 12'sd1138, 11'sd1016}},
{{12'sd1216, 8'sd71, 11'sd-779}, {12'sd-1893, 13'sd2083, 12'sd-1880}, {12'sd-1400, 12'sd1873, 12'sd-1468}},
{{9'sd-185, 13'sd-3270, 12'sd-1646}, {12'sd-1157, 12'sd-1442, 13'sd-2427}, {12'sd1524, 8'sd-85, 13'sd2385}},
{{13'sd-2374, 13'sd3283, 13'sd-3347}, {13'sd-2445, 13'sd2895, 12'sd1359}, {11'sd725, 12'sd1187, 12'sd-1055}},
{{11'sd887, 13'sd2638, 9'sd214}, {12'sd-1559, 13'sd2623, 13'sd-2954}, {13'sd-2109, 12'sd1272, 10'sd449}}},
{
{{11'sd-914, 12'sd1334, 9'sd230}, {11'sd-777, 12'sd1497, 12'sd-1889}, {12'sd-1644, 10'sd-509, 13'sd-2523}},
{{13'sd2863, 13'sd-2398, 8'sd-72}, {12'sd-1277, 9'sd-176, 12'sd-1064}, {12'sd1699, 13'sd-2671, 10'sd297}},
{{13'sd2097, 12'sd1378, 13'sd-2356}, {12'sd1492, 12'sd-1080, 13'sd-2256}, {7'sd40, 12'sd-1548, 11'sd-950}},
{{12'sd1883, 11'sd-772, 12'sd-1628}, {10'sd-415, 12'sd-1514, 9'sd-253}, {12'sd1839, 10'sd-295, 13'sd2791}},
{{13'sd-3062, 12'sd-1196, 11'sd1021}, {14'sd-5208, 9'sd-241, 13'sd-3115}, {13'sd-2438, 10'sd472, 14'sd-4277}},
{{12'sd1298, 12'sd-1757, 11'sd-912}, {13'sd-2550, 12'sd1246, 8'sd118}, {12'sd1105, 10'sd-260, 12'sd-1451}},
{{12'sd1531, 12'sd1816, 12'sd1564}, {11'sd556, 11'sd960, 10'sd-500}, {12'sd1144, 14'sd4199, 13'sd3001}},
{{11'sd584, 12'sd1501, 12'sd1554}, {12'sd-1290, 7'sd32, 12'sd1401}, {13'sd2707, 10'sd-451, 9'sd-129}},
{{10'sd270, 12'sd-1994, 13'sd-2174}, {13'sd-2098, 12'sd-1369, 12'sd1081}, {12'sd-1629, 12'sd-1172, 11'sd636}},
{{9'sd-184, 8'sd76, 9'sd238}, {12'sd-1994, 12'sd1150, 13'sd2266}, {12'sd-1024, 10'sd-364, 13'sd-2206}},
{{13'sd3021, 12'sd1236, 12'sd1511}, {9'sd250, 12'sd1219, 11'sd652}, {13'sd2098, 13'sd2472, 12'sd1965}},
{{13'sd2778, 12'sd-1809, 13'sd2099}, {12'sd-1394, 13'sd-2682, 12'sd1631}, {11'sd791, 10'sd338, 9'sd-136}},
{{13'sd-3167, 12'sd1354, 11'sd-550}, {11'sd936, 13'sd-3176, 12'sd-2039}, {10'sd-386, 13'sd-2661, 10'sd388}},
{{8'sd-87, 11'sd-649, 13'sd2663}, {13'sd2309, 10'sd-416, 12'sd1253}, {13'sd-2183, 12'sd-1460, 13'sd2227}},
{{14'sd-4266, 9'sd-233, 12'sd1683}, {13'sd-3156, 13'sd2300, 11'sd-718}, {13'sd-2495, 11'sd-761, 11'sd-564}},
{{10'sd-268, 12'sd-1732, 11'sd-900}, {11'sd-550, 12'sd1378, 12'sd-1220}, {11'sd-876, 11'sd888, 6'sd-17}},
{{13'sd2896, 11'sd662, 13'sd-2458}, {13'sd2515, 12'sd-1288, 13'sd2567}, {13'sd2424, 13'sd2234, 10'sd-312}},
{{13'sd-2453, 10'sd-455, 12'sd-1721}, {13'sd-2868, 12'sd-1464, 13'sd-2400}, {13'sd-2997, 12'sd1832, 12'sd-1622}},
{{8'sd124, 11'sd-801, 10'sd-498}, {12'sd-1458, 13'sd2930, 11'sd640}, {12'sd-1468, 13'sd2744, 12'sd1128}},
{{13'sd-2408, 13'sd-2113, 9'sd-174}, {9'sd-148, 13'sd2189, 12'sd-1879}, {11'sd-658, 12'sd1078, 13'sd-2058}},
{{8'sd109, 10'sd-341, 10'sd359}, {13'sd-2799, 13'sd-2120, 10'sd-481}, {12'sd-1494, 13'sd2823, 13'sd-2116}},
{{10'sd-444, 13'sd-2622, 10'sd338}, {11'sd855, 10'sd442, 12'sd-1529}, {12'sd-1915, 13'sd2665, 13'sd-2355}},
{{12'sd-1729, 9'sd150, 12'sd-1508}, {11'sd597, 12'sd-1075, 11'sd-753}, {12'sd2046, 13'sd-2822, 12'sd-1568}},
{{12'sd1197, 13'sd2345, 12'sd2012}, {12'sd1791, 12'sd-1251, 11'sd854}, {12'sd1903, 12'sd-1957, 10'sd-362}},
{{10'sd471, 12'sd-1623, 10'sd306}, {12'sd-1917, 13'sd2156, 12'sd-1756}, {12'sd-2041, 12'sd-1961, 10'sd-402}},
{{12'sd1506, 11'sd-733, 13'sd-2417}, {12'sd-1806, 13'sd-2394, 11'sd-690}, {11'sd852, 11'sd826, 11'sd722}},
{{13'sd2271, 11'sd831, 13'sd3586}, {12'sd-1830, 12'sd1111, 11'sd-828}, {12'sd1135, 11'sd-689, 11'sd933}},
{{9'sd173, 13'sd2443, 12'sd-1171}, {13'sd-2178, 10'sd-363, 12'sd1533}, {4'sd-7, 12'sd-1484, 8'sd90}},
{{12'sd1496, 11'sd-564, 13'sd2611}, {13'sd2507, 13'sd3306, 11'sd736}, {13'sd2141, 13'sd2171, 9'sd142}},
{{11'sd708, 12'sd1579, 11'sd-889}, {7'sd-49, 13'sd2670, 11'sd1003}, {13'sd2108, 13'sd2333, 12'sd1410}},
{{12'sd-1848, 13'sd-2416, 12'sd-1577}, {12'sd1712, 13'sd2450, 12'sd1869}, {13'sd-2284, 13'sd2454, 12'sd2030}},
{{12'sd-1937, 11'sd663, 12'sd-1175}, {13'sd2853, 13'sd2635, 3'sd-3}, {12'sd2016, 13'sd2750, 12'sd-1284}},
{{8'sd-124, 13'sd2063, 12'sd1457}, {13'sd-2450, 12'sd-1450, 10'sd-460}, {7'sd-56, 12'sd-1705, 11'sd-828}},
{{12'sd-1441, 12'sd-1348, 12'sd2007}, {10'sd349, 12'sd1348, 10'sd305}, {11'sd-651, 12'sd-1583, 12'sd1622}},
{{13'sd2323, 11'sd-734, 9'sd-184}, {11'sd-780, 12'sd1622, 13'sd3099}, {10'sd412, 8'sd100, 11'sd-516}},
{{12'sd-1286, 10'sd-280, 13'sd2668}, {12'sd-1162, 13'sd2835, 12'sd1888}, {8'sd-92, 12'sd1812, 12'sd1545}},
{{11'sd-768, 11'sd-690, 11'sd514}, {8'sd-74, 13'sd2210, 12'sd1470}, {12'sd-1941, 13'sd2840, 10'sd-369}},
{{13'sd-2700, 12'sd1550, 11'sd-540}, {12'sd1862, 12'sd-1274, 12'sd-1486}, {12'sd-1918, 13'sd-2856, 12'sd-1918}},
{{13'sd2255, 12'sd1330, 12'sd-1165}, {12'sd-1503, 9'sd197, 13'sd2375}, {12'sd-1203, 13'sd2316, 9'sd-130}},
{{12'sd-1631, 13'sd-2897, 12'sd1662}, {12'sd-1967, 11'sd607, 9'sd241}, {13'sd2062, 10'sd307, 12'sd1246}},
{{11'sd-873, 13'sd-3122, 13'sd-2679}, {10'sd-373, 11'sd796, 11'sd-988}, {13'sd2402, 12'sd1109, 12'sd1231}},
{{12'sd-1671, 12'sd-2025, 12'sd-1414}, {9'sd-223, 12'sd-1614, 13'sd-2261}, {12'sd-1042, 12'sd1743, 12'sd-1982}},
{{10'sd-381, 12'sd1906, 12'sd-1373}, {12'sd-1630, 8'sd78, 9'sd-212}, {12'sd1647, 11'sd690, 13'sd2555}},
{{11'sd907, 11'sd729, 13'sd3949}, {12'sd-1563, 12'sd1500, 12'sd1473}, {9'sd-133, 9'sd-228, 13'sd-2163}},
{{13'sd2227, 12'sd-1059, 13'sd2368}, {9'sd-224, 12'sd1671, 12'sd1657}, {11'sd-991, 9'sd221, 9'sd155}},
{{12'sd1921, 11'sd-751, 12'sd1598}, {12'sd1958, 12'sd1188, 13'sd-2529}, {12'sd-1448, 10'sd401, 7'sd-61}},
{{11'sd650, 12'sd-1829, 11'sd715}, {12'sd1134, 6'sd26, 11'sd524}, {11'sd-624, 12'sd1781, 11'sd-811}},
{{11'sd-1006, 11'sd-708, 13'sd2789}, {12'sd1133, 13'sd-2440, 11'sd1022}, {11'sd-567, 11'sd-835, 12'sd-1422}},
{{10'sd392, 13'sd2269, 10'sd-361}, {11'sd938, 12'sd1987, 11'sd-625}, {11'sd752, 11'sd-821, 11'sd822}},
{{13'sd-2136, 12'sd1208, 12'sd-1364}, {11'sd533, 12'sd-1222, 13'sd2663}, {13'sd-3098, 13'sd2559, 7'sd-63}},
{{12'sd1691, 13'sd2482, 12'sd1673}, {9'sd232, 12'sd-1611, 13'sd2369}, {11'sd-533, 11'sd648, 13'sd2434}},
{{11'sd-649, 11'sd-926, 13'sd-2115}, {12'sd1357, 13'sd-2150, 12'sd-1261}, {13'sd2728, 12'sd-1115, 13'sd2236}},
{{12'sd-1908, 11'sd-944, 13'sd-2306}, {9'sd-221, 12'sd1194, 11'sd-1002}, {7'sd47, 12'sd-1960, 12'sd1969}},
{{9'sd-146, 12'sd1706, 13'sd2436}, {12'sd1881, 13'sd2697, 12'sd-1125}, {12'sd1572, 12'sd1430, 12'sd1601}},
{{14'sd-4676, 9'sd248, 12'sd-1732}, {11'sd-873, 12'sd1157, 13'sd-2152}, {11'sd633, 13'sd3330, 13'sd-2493}},
{{13'sd2549, 9'sd-214, 11'sd991}, {10'sd278, 13'sd2904, 13'sd2086}, {4'sd5, 10'sd431, 10'sd424}},
{{8'sd119, 14'sd-4396, 14'sd-4324}, {10'sd339, 13'sd-3253, 13'sd-3625}, {12'sd-1385, 12'sd-1600, 10'sd-374}},
{{12'sd2027, 12'sd1408, 12'sd-1285}, {11'sd-977, 13'sd-2210, 13'sd-3105}, {12'sd1435, 12'sd-1662, 10'sd-443}},
{{13'sd2206, 12'sd1236, 11'sd-819}, {12'sd1588, 13'sd-2123, 13'sd-2395}, {12'sd-1893, 13'sd-2546, 11'sd576}},
{{13'sd-2672, 11'sd841, 11'sd-728}, {12'sd-2010, 13'sd3358, 9'sd144}, {12'sd1870, 13'sd2549, 12'sd-1425}},
{{12'sd-1316, 12'sd-1576, 11'sd-544}, {13'sd-2052, 9'sd-250, 13'sd-2298}, {11'sd-849, 13'sd-2473, 12'sd-1899}},
{{10'sd-413, 13'sd-2963, 12'sd-1210}, {9'sd-237, 10'sd416, 12'sd1698}, {12'sd-1389, 12'sd1415, 13'sd-2061}},
{{12'sd-1996, 12'sd1830, 12'sd-1211}, {13'sd-2165, 11'sd-632, 12'sd1818}, {12'sd1670, 12'sd-1166, 9'sd131}},
{{12'sd-1477, 13'sd3495, 12'sd-1588}, {10'sd428, 8'sd67, 10'sd336}, {11'sd-829, 12'sd1663, 13'sd2902}}},
{
{{12'sd1717, 13'sd-2315, 12'sd-1122}, {10'sd-351, 12'sd1654, 13'sd-2671}, {12'sd-1417, 11'sd-1013, 9'sd227}},
{{12'sd-1389, 10'sd484, 13'sd-2481}, {13'sd-2113, 12'sd1833, 12'sd1787}, {12'sd1183, 13'sd2334, 13'sd-2717}},
{{13'sd-2187, 13'sd-2257, 12'sd-1570}, {12'sd1542, 13'sd-2654, 12'sd1927}, {12'sd1927, 11'sd-770, 12'sd1868}},
{{9'sd-239, 9'sd-163, 13'sd2512}, {12'sd1943, 12'sd-1866, 12'sd-1312}, {12'sd-1582, 12'sd-1547, 12'sd-1621}},
{{10'sd302, 12'sd-1995, 12'sd1231}, {13'sd-3532, 13'sd-4062, 12'sd-1088}, {13'sd-2272, 12'sd-1855, 12'sd-1170}},
{{12'sd-1416, 10'sd-472, 13'sd3139}, {13'sd-4021, 12'sd1139, 12'sd-1330}, {12'sd-1506, 12'sd-1274, 13'sd-2424}},
{{13'sd-2380, 10'sd459, 13'sd2910}, {12'sd-1658, 12'sd1307, 11'sd-845}, {12'sd-1499, 12'sd1075, 11'sd-794}},
{{10'sd415, 13'sd-2403, 12'sd1329}, {13'sd2393, 11'sd1013, 11'sd914}, {12'sd1104, 12'sd-1595, 12'sd-1147}},
{{11'sd-650, 12'sd1118, 12'sd-2034}, {11'sd-657, 13'sd2137, 13'sd2370}, {12'sd-1376, 10'sd425, 12'sd1942}},
{{12'sd-1844, 11'sd620, 12'sd1240}, {13'sd2223, 13'sd2193, 13'sd-2886}, {13'sd2370, 13'sd-2327, 12'sd1067}},
{{13'sd2101, 12'sd1710, 9'sd-162}, {13'sd2109, 13'sd-2459, 9'sd175}, {13'sd3509, 11'sd868, 13'sd2146}},
{{11'sd-898, 12'sd1849, 11'sd-767}, {9'sd-131, 13'sd-2539, 12'sd1411}, {8'sd111, 12'sd-1874, 12'sd1131}},
{{12'sd-1177, 5'sd9, 11'sd-714}, {12'sd-1222, 13'sd-2859, 12'sd1519}, {12'sd1833, 11'sd523, 13'sd-2761}},
{{12'sd1745, 12'sd1713, 12'sd1280}, {12'sd1424, 12'sd1235, 12'sd-1323}, {12'sd1260, 13'sd2320, 12'sd-1743}},
{{9'sd-198, 11'sd-734, 13'sd2055}, {11'sd-844, 12'sd-1978, 13'sd2050}, {13'sd-3010, 12'sd1233, 11'sd725}},
{{10'sd408, 12'sd1644, 10'sd-310}, {10'sd274, 12'sd1975, 10'sd305}, {10'sd-368, 8'sd-110, 13'sd-2594}},
{{13'sd2299, 13'sd3038, 11'sd974}, {12'sd-1269, 12'sd-1992, 10'sd353}, {11'sd603, 11'sd800, 11'sd-796}},
{{13'sd-2839, 12'sd1770, 12'sd1973}, {10'sd-286, 13'sd-3416, 12'sd-1954}, {13'sd-3491, 12'sd-1094, 12'sd1866}},
{{11'sd-686, 13'sd2521, 12'sd-2045}, {12'sd1333, 12'sd-1032, 10'sd-437}, {12'sd1871, 10'sd313, 8'sd100}},
{{11'sd814, 13'sd2653, 10'sd-268}, {13'sd-2284, 12'sd1567, 13'sd-2577}, {12'sd-1356, 10'sd-502, 13'sd-2693}},
{{10'sd349, 12'sd-2045, 12'sd-1623}, {11'sd933, 10'sd-275, 12'sd1520}, {9'sd-191, 13'sd-2203, 12'sd1692}},
{{13'sd2437, 12'sd-1231, 10'sd366}, {13'sd-2466, 11'sd-963, 11'sd630}, {9'sd-188, 2'sd1, 12'sd-2045}},
{{6'sd-29, 11'sd933, 13'sd-2474}, {13'sd2312, 13'sd-2554, 12'sd1108}, {12'sd-1452, 12'sd1499, 13'sd-2235}},
{{10'sd-454, 12'sd-1498, 13'sd-2130}, {9'sd-251, 13'sd2122, 12'sd1186}, {12'sd-1234, 9'sd137, 11'sd-1014}},
{{10'sd301, 13'sd2311, 10'sd-494}, {12'sd1322, 5'sd-10, 11'sd-641}, {11'sd729, 12'sd-1401, 13'sd-2847}},
{{13'sd2229, 12'sd-1930, 12'sd-1894}, {12'sd-1230, 12'sd1278, 11'sd624}, {13'sd2271, 13'sd-2338, 11'sd-693}},
{{13'sd2982, 12'sd-2019, 13'sd2625}, {12'sd-1265, 10'sd272, 11'sd-593}, {12'sd1062, 13'sd3700, 13'sd2484}},
{{12'sd-1094, 11'sd612, 9'sd-216}, {13'sd-2287, 12'sd-1683, 13'sd-2886}, {13'sd-2321, 13'sd-2238, 12'sd1335}},
{{9'sd-131, 13'sd2952, 11'sd874}, {13'sd-2063, 12'sd1046, 13'sd-2157}, {12'sd-1318, 13'sd2137, 11'sd-975}},
{{12'sd1527, 12'sd-1455, 13'sd-3451}, {11'sd975, 12'sd-1631, 10'sd298}, {13'sd2456, 8'sd98, 13'sd2656}},
{{13'sd-2086, 13'sd2864, 12'sd-1506}, {8'sd-71, 9'sd236, 12'sd1921}, {11'sd821, 12'sd1735, 11'sd-871}},
{{13'sd3212, 13'sd2049, 13'sd2751}, {11'sd-637, 13'sd2097, 8'sd115}, {9'sd208, 12'sd1604, 12'sd1271}},
{{13'sd-2121, 9'sd148, 11'sd656}, {12'sd2001, 12'sd-1704, 12'sd-1989}, {12'sd-1599, 10'sd-380, 11'sd951}},
{{10'sd-355, 13'sd2246, 11'sd-543}, {12'sd-1828, 12'sd-1078, 9'sd178}, {12'sd-1244, 12'sd-1435, 13'sd-2588}},
{{13'sd2259, 11'sd591, 10'sd-407}, {13'sd-2445, 12'sd-1743, 11'sd-1012}, {13'sd-2563, 12'sd-1914, 11'sd-829}},
{{12'sd1954, 12'sd-1059, 12'sd2012}, {13'sd-2470, 11'sd-514, 12'sd-1938}, {13'sd-2759, 10'sd-265, 12'sd1798}},
{{10'sd-276, 13'sd3230, 13'sd2265}, {6'sd23, 10'sd449, 8'sd-118}, {12'sd-1530, 8'sd-99, 13'sd3016}},
{{12'sd-1542, 10'sd265, 13'sd-2227}, {13'sd-3251, 11'sd-625, 12'sd-1346}, {12'sd1902, 13'sd-2410, 13'sd-2805}},
{{12'sd1106, 11'sd-679, 11'sd875}, {12'sd-1091, 12'sd-1103, 10'sd488}, {12'sd-1787, 9'sd204, 12'sd-1801}},
{{13'sd-2650, 12'sd-1941, 13'sd-2459}, {12'sd-1732, 12'sd-1919, 12'sd-1689}, {13'sd2832, 11'sd554, 13'sd-2370}},
{{12'sd-1432, 12'sd-1415, 12'sd1464}, {12'sd-1195, 11'sd602, 13'sd-2308}, {13'sd-3299, 10'sd448, 13'sd-3130}},
{{12'sd1458, 13'sd2669, 12'sd1294}, {12'sd1373, 12'sd-1740, 9'sd-193}, {10'sd462, 9'sd211, 10'sd278}},
{{11'sd-905, 10'sd-501, 10'sd-335}, {12'sd1787, 10'sd-364, 11'sd-925}, {13'sd2196, 12'sd1065, 11'sd-642}},
{{13'sd3722, 13'sd3946, 14'sd4755}, {13'sd3618, 13'sd3063, 7'sd45}, {14'sd7232, 14'sd6091, 14'sd4422}},
{{10'sd-505, 10'sd331, 8'sd-68}, {12'sd-1256, 13'sd-2280, 13'sd2102}, {13'sd2339, 12'sd2043, 13'sd-2624}},
{{12'sd1393, 13'sd2408, 9'sd218}, {11'sd574, 12'sd1450, 12'sd1561}, {13'sd2057, 9'sd-138, 12'sd-1590}},
{{10'sd-269, 12'sd-1563, 12'sd-1536}, {13'sd2345, 10'sd-455, 13'sd-2201}, {11'sd660, 11'sd812, 11'sd-890}},
{{12'sd1137, 13'sd2138, 8'sd98}, {13'sd-3500, 12'sd1123, 9'sd223}, {13'sd-3152, 13'sd2143, 12'sd-1639}},
{{12'sd-1435, 11'sd-546, 13'sd2547}, {11'sd937, 11'sd-845, 13'sd2721}, {11'sd686, 12'sd1259, 11'sd688}},
{{10'sd-288, 13'sd-2522, 12'sd1247}, {13'sd2251, 13'sd3338, 12'sd-1118}, {12'sd-1669, 12'sd1779, 13'sd-2816}},
{{13'sd2473, 13'sd-2442, 13'sd2258}, {12'sd1315, 12'sd-1781, 12'sd1339}, {12'sd1792, 13'sd2430, 13'sd-2715}},
{{12'sd-1992, 12'sd2044, 10'sd-411}, {10'sd-397, 10'sd377, 13'sd2699}, {11'sd-701, 13'sd2502, 12'sd-1816}},
{{13'sd2270, 12'sd1839, 10'sd-281}, {12'sd-1494, 12'sd1191, 13'sd-2820}, {13'sd3290, 11'sd-976, 12'sd-1715}},
{{13'sd-2444, 13'sd2720, 13'sd2064}, {13'sd2569, 10'sd442, 11'sd-937}, {11'sd542, 13'sd-2291, 12'sd-1777}},
{{12'sd-1554, 12'sd1489, 13'sd-3224}, {9'sd254, 12'sd-1202, 13'sd-3589}, {13'sd-4069, 12'sd1294, 13'sd-3063}},
{{12'sd1063, 10'sd405, 8'sd-112}, {12'sd-1237, 11'sd925, 11'sd-670}, {12'sd-1801, 12'sd1540, 12'sd-1703}},
{{11'sd-939, 9'sd171, 8'sd121}, {12'sd1069, 8'sd85, 13'sd-2208}, {12'sd1962, 11'sd772, 11'sd911}},
{{12'sd-1347, 11'sd654, 12'sd1610}, {10'sd-369, 12'sd-1900, 12'sd-1864}, {11'sd760, 13'sd-2938, 11'sd-729}},
{{12'sd-1779, 12'sd1189, 8'sd-105}, {12'sd-1343, 11'sd857, 13'sd-2714}, {10'sd-420, 12'sd-1659, 13'sd2611}},
{{13'sd-2461, 13'sd2452, 12'sd-1271}, {13'sd-2095, 10'sd404, 13'sd2221}, {14'sd-4395, 13'sd-3851, 12'sd1133}},
{{12'sd1134, 12'sd-1995, 12'sd-1475}, {13'sd-2088, 11'sd719, 12'sd1285}, {10'sd413, 12'sd-1054, 10'sd-286}},
{{13'sd-2054, 10'sd-344, 13'sd-2652}, {11'sd-894, 13'sd-2465, 11'sd-642}, {12'sd2041, 12'sd-1529, 12'sd1674}},
{{13'sd2130, 12'sd-1941, 13'sd2357}, {11'sd-744, 12'sd-1451, 12'sd-1774}, {13'sd-2565, 13'sd-2850, 12'sd-1552}},
{{13'sd3086, 10'sd262, 12'sd1966}, {13'sd2859, 12'sd2023, 12'sd1926}, {13'sd3042, 7'sd55, 13'sd2200}}},
{
{{12'sd1281, 13'sd2690, 13'sd-2781}, {12'sd1378, 12'sd1304, 13'sd-2230}, {13'sd2215, 11'sd-695, 12'sd-1202}},
{{13'sd3265, 13'sd2867, 13'sd3146}, {12'sd1315, 12'sd-1781, 11'sd1017}, {12'sd-1290, 8'sd126, 13'sd-2660}},
{{12'sd-1374, 12'sd1358, 13'sd-2084}, {12'sd-1452, 11'sd-632, 12'sd1400}, {13'sd2372, 13'sd-2092, 12'sd1165}},
{{13'sd2290, 12'sd-1486, 11'sd-687}, {12'sd-1407, 11'sd-762, 12'sd-1162}, {10'sd416, 10'sd-351, 12'sd-1407}},
{{11'sd781, 13'sd2558, 10'sd411}, {13'sd2808, 13'sd3583, 12'sd1684}, {10'sd342, 10'sd-273, 11'sd632}},
{{10'sd-470, 12'sd-1632, 11'sd666}, {13'sd3474, 12'sd-1728, 13'sd2369}, {12'sd-1675, 12'sd1125, 12'sd1680}},
{{11'sd-942, 10'sd-276, 12'sd1555}, {11'sd948, 12'sd2004, 12'sd-1335}, {11'sd-692, 14'sd-4956, 14'sd-4099}},
{{11'sd933, 11'sd-601, 10'sd277}, {11'sd731, 12'sd-1695, 12'sd1575}, {12'sd-1244, 12'sd1496, 13'sd-2147}},
{{13'sd2311, 11'sd-911, 5'sd-12}, {10'sd-349, 11'sd631, 13'sd-2347}, {12'sd-1725, 12'sd-1199, 12'sd-1408}},
{{13'sd-2761, 8'sd-76, 12'sd1896}, {11'sd977, 12'sd1449, 12'sd-1924}, {13'sd-2616, 12'sd-1346, 9'sd-223}},
{{11'sd769, 13'sd2674, 12'sd1631}, {10'sd476, 13'sd2946, 13'sd-3013}, {12'sd1163, 12'sd-1312, 13'sd-3500}},
{{11'sd811, 12'sd1895, 11'sd-738}, {9'sd-242, 13'sd2845, 13'sd2623}, {13'sd3012, 13'sd3135, 11'sd-983}},
{{11'sd758, 13'sd3522, 11'sd-834}, {12'sd-1175, 12'sd-1492, 12'sd-1094}, {12'sd-1912, 13'sd-3079, 11'sd573}},
{{11'sd609, 12'sd-1768, 13'sd2303}, {9'sd-232, 8'sd94, 10'sd-314}, {11'sd646, 13'sd2939, 8'sd115}},
{{13'sd4081, 6'sd20, 11'sd-834}, {7'sd-63, 12'sd1204, 10'sd507}, {10'sd492, 11'sd521, 11'sd-763}},
{{13'sd-3355, 12'sd1237, 11'sd-599}, {13'sd3438, 6'sd-22, 12'sd1492}, {8'sd-66, 11'sd779, 11'sd-561}},
{{12'sd-1842, 11'sd-715, 10'sd-371}, {12'sd1917, 12'sd1254, 13'sd2947}, {12'sd-1156, 13'sd3097, 13'sd2789}},
{{6'sd-28, 12'sd1615, 12'sd1802}, {13'sd2395, 13'sd2292, 11'sd523}, {11'sd-546, 12'sd-1516, 8'sd-68}},
{{10'sd457, 13'sd-2378, 11'sd732}, {13'sd-2648, 12'sd1654, 9'sd185}, {13'sd-2578, 10'sd-296, 11'sd648}},
{{13'sd-2425, 13'sd-2407, 11'sd-545}, {13'sd-2707, 9'sd-189, 11'sd690}, {12'sd1436, 12'sd-1652, 9'sd195}},
{{12'sd-1101, 11'sd941, 12'sd-1433}, {12'sd1198, 9'sd173, 12'sd-1162}, {10'sd-437, 13'sd-2720, 13'sd-2529}},
{{12'sd1471, 11'sd-873, 9'sd-145}, {12'sd1924, 11'sd928, 12'sd-1794}, {13'sd2796, 13'sd2997, 13'sd3262}},
{{10'sd465, 13'sd-2146, 11'sd-633}, {11'sd-879, 12'sd-1864, 11'sd-534}, {13'sd2702, 12'sd1673, 12'sd1213}},
{{10'sd-391, 13'sd-2679, 9'sd-165}, {13'sd-2293, 3'sd-3, 11'sd661}, {11'sd684, 12'sd1190, 12'sd1582}},
{{12'sd-1768, 10'sd371, 11'sd-727}, {12'sd-1279, 11'sd518, 12'sd1696}, {12'sd1535, 13'sd-2523, 10'sd381}},
{{12'sd1766, 13'sd2117, 12'sd-1523}, {10'sd-418, 12'sd1232, 12'sd1357}, {12'sd-1711, 11'sd854, 13'sd-2845}},
{{13'sd2651, 13'sd-2301, 12'sd1413}, {12'sd1764, 13'sd-3538, 12'sd-1411}, {12'sd-1687, 12'sd-1952, 13'sd-2735}},
{{12'sd-1815, 12'sd1756, 11'sd-898}, {13'sd2654, 13'sd3196, 12'sd-1555}, {12'sd-1277, 12'sd-1089, 13'sd-2345}},
{{13'sd2182, 11'sd993, 13'sd2120}, {12'sd-1065, 13'sd-2413, 8'sd-66}, {12'sd1782, 12'sd1425, 10'sd357}},
{{12'sd-1260, 13'sd2318, 7'sd-42}, {12'sd-1945, 13'sd2386, 12'sd1259}, {13'sd-3786, 12'sd1105, 6'sd-29}},
{{13'sd-3013, 10'sd313, 12'sd-1116}, {13'sd-2112, 13'sd-2531, 11'sd-940}, {10'sd-439, 11'sd-961, 13'sd2290}},
{{12'sd1822, 12'sd1326, 13'sd2828}, {12'sd1880, 12'sd-1872, 12'sd-1413}, {12'sd-1149, 11'sd-525, 13'sd-2456}},
{{13'sd-2061, 13'sd-2200, 12'sd1091}, {5'sd11, 12'sd1300, 10'sd276}, {11'sd609, 12'sd1728, 11'sd-540}},
{{12'sd-1440, 12'sd-1174, 13'sd-2753}, {9'sd170, 12'sd1638, 12'sd1418}, {11'sd-884, 12'sd1569, 11'sd749}},
{{13'sd-3312, 10'sd408, 12'sd1052}, {9'sd192, 12'sd1605, 11'sd-789}, {11'sd-524, 9'sd214, 14'sd4184}},
{{11'sd578, 12'sd-1259, 11'sd739}, {9'sd213, 11'sd824, 9'sd-192}, {12'sd1453, 12'sd1476, 10'sd-312}},
{{12'sd1224, 12'sd-2028, 13'sd-2233}, {13'sd-2335, 12'sd-1486, 12'sd-1317}, {12'sd-1608, 10'sd256, 12'sd-2038}},
{{11'sd-781, 13'sd-2918, 12'sd-1593}, {12'sd1640, 9'sd-237, 12'sd-1283}, {12'sd1499, 12'sd1424, 12'sd1420}},
{{11'sd-585, 9'sd-144, 10'sd-377}, {13'sd2249, 12'sd-1783, 12'sd-1524}, {11'sd975, 12'sd-1247, 11'sd834}},
{{12'sd1956, 13'sd2094, 13'sd2514}, {12'sd-1608, 11'sd526, 10'sd-504}, {13'sd-2656, 11'sd-598, 12'sd-1863}},
{{10'sd388, 12'sd1167, 11'sd-571}, {10'sd-406, 10'sd411, 11'sd-707}, {12'sd1318, 13'sd-3161, 10'sd356}},
{{11'sd-969, 13'sd3592, 7'sd47}, {11'sd792, 12'sd1531, 10'sd356}, {11'sd749, 12'sd-1990, 13'sd-2532}},
{{12'sd-1863, 10'sd-340, 10'sd-293}, {11'sd569, 12'sd-1289, 13'sd-2581}, {10'sd459, 13'sd-2497, 13'sd-3442}},
{{14'sd7427, 13'sd4084, 9'sd-253}, {14'sd5406, 11'sd905, 12'sd1928}, {13'sd3967, 13'sd2371, 13'sd3107}},
{{12'sd-1467, 11'sd915, 11'sd632}, {12'sd-1458, 7'sd-57, 13'sd2650}, {12'sd-2020, 12'sd1092, 12'sd1213}},
{{10'sd-387, 12'sd-1507, 11'sd623}, {11'sd668, 11'sd837, 5'sd10}, {12'sd-1379, 12'sd-1911, 13'sd3560}},
{{13'sd2327, 9'sd162, 13'sd-2909}, {13'sd2477, 12'sd-1739, 13'sd2638}, {13'sd-3285, 11'sd-939, 10'sd344}},
{{13'sd2325, 13'sd-2357, 12'sd1800}, {13'sd-2068, 13'sd2754, 12'sd1827}, {13'sd2352, 12'sd1428, 11'sd-682}},
{{13'sd-2080, 11'sd-1016, 12'sd-1774}, {13'sd-2484, 11'sd-632, 10'sd272}, {13'sd-2489, 13'sd-2881, 13'sd-3071}},
{{11'sd870, 13'sd-2223, 11'sd915}, {11'sd736, 11'sd870, 11'sd673}, {13'sd2294, 11'sd-638, 13'sd2309}},
{{11'sd846, 13'sd-3212, 13'sd-2250}, {11'sd938, 10'sd481, 12'sd2047}, {12'sd-1139, 11'sd771, 13'sd3305}},
{{10'sd488, 12'sd1906, 13'sd-2363}, {10'sd326, 12'sd-1092, 12'sd-1181}, {10'sd-502, 12'sd1670, 12'sd-1084}},
{{11'sd1022, 11'sd-820, 10'sd-324}, {13'sd-3321, 13'sd2361, 12'sd-1208}, {9'sd-186, 12'sd-1357, 12'sd1580}},
{{12'sd1958, 10'sd-303, 13'sd2884}, {13'sd2150, 13'sd-2325, 13'sd2129}, {12'sd1230, 13'sd-2262, 13'sd2491}},
{{12'sd1980, 11'sd777, 12'sd-1695}, {12'sd1113, 11'sd734, 10'sd388}, {13'sd-2423, 13'sd-2546, 14'sd-4734}},
{{12'sd-1870, 10'sd-258, 11'sd-905}, {13'sd-2322, 10'sd-297, 9'sd176}, {12'sd1060, 12'sd1119, 12'sd-1713}},
{{10'sd-410, 12'sd1949, 11'sd1021}, {9'sd148, 11'sd-722, 13'sd3487}, {12'sd-1394, 11'sd884, 13'sd2965}},
{{11'sd-980, 13'sd2858, 12'sd2037}, {13'sd3584, 10'sd-416, 13'sd3100}, {10'sd-431, 12'sd-1422, 13'sd2579}},
{{13'sd2836, 11'sd877, 11'sd-514}, {13'sd2471, 11'sd-594, 12'sd1226}, {11'sd561, 13'sd-2115, 10'sd-408}},
{{12'sd1690, 13'sd-2160, 12'sd-1255}, {11'sd793, 10'sd401, 11'sd519}, {14'sd-5044, 12'sd-1038, 14'sd-4481}},
{{12'sd1028, 11'sd659, 12'sd1246}, {11'sd-590, 12'sd-1200, 12'sd-1680}, {12'sd1231, 11'sd-548, 13'sd3186}},
{{11'sd945, 13'sd-2094, 13'sd-2683}, {12'sd1953, 11'sd865, 13'sd-2572}, {9'sd-243, 11'sd-629, 11'sd547}},
{{13'sd2786, 13'sd-2359, 12'sd-1026}, {12'sd1052, 11'sd-959, 13'sd2392}, {12'sd1027, 13'sd-2159, 11'sd-675}},
{{12'sd-1953, 12'sd2030, 11'sd-779}, {10'sd284, 11'sd839, 11'sd-693}, {11'sd717, 10'sd272, 13'sd-2333}}},
{
{{12'sd-1214, 10'sd-480, 13'sd2884}, {10'sd-499, 13'sd-2790, 12'sd-1813}, {12'sd1241, 12'sd1237, 10'sd319}},
{{12'sd-2014, 10'sd286, 12'sd-1375}, {13'sd-2390, 13'sd-2268, 12'sd1513}, {12'sd1694, 13'sd-2632, 12'sd-1032}},
{{13'sd3072, 7'sd49, 12'sd-1050}, {11'sd927, 12'sd1370, 12'sd-1760}, {11'sd522, 13'sd2299, 12'sd-1239}},
{{10'sd-362, 12'sd1546, 12'sd-1322}, {12'sd1474, 11'sd-933, 12'sd-1037}, {12'sd-1071, 12'sd1867, 11'sd1021}},
{{13'sd-3534, 12'sd-1289, 11'sd-543}, {13'sd-2332, 13'sd-2395, 10'sd-260}, {5'sd15, 13'sd-2578, 13'sd-3242}},
{{12'sd1291, 12'sd1267, 12'sd-1173}, {13'sd-2726, 12'sd-1902, 12'sd-1563}, {12'sd-2001, 8'sd-112, 12'sd1038}},
{{13'sd-3822, 13'sd-3174, 10'sd400}, {12'sd1284, 11'sd885, 13'sd2319}, {12'sd1906, 12'sd1990, 13'sd2571}},
{{12'sd-2002, 11'sd-906, 12'sd1741}, {12'sd-1559, 11'sd950, 11'sd842}, {11'sd892, 12'sd-1602, 12'sd1348}},
{{12'sd-1097, 11'sd-1006, 13'sd2293}, {13'sd-2318, 13'sd-2180, 13'sd-2419}, {12'sd1255, 11'sd588, 9'sd208}},
{{12'sd1324, 11'sd-985, 12'sd1560}, {12'sd-1178, 12'sd-1282, 12'sd1211}, {5'sd-14, 13'sd-2462, 10'sd-327}},
{{11'sd761, 13'sd-2328, 8'sd-93}, {11'sd515, 10'sd-259, 10'sd386}, {12'sd-1202, 12'sd-2039, 13'sd2132}},
{{13'sd2991, 11'sd850, 13'sd2188}, {12'sd1027, 12'sd-1926, 7'sd-55}, {13'sd-2442, 13'sd2515, 13'sd-2120}},
{{12'sd-1893, 11'sd-748, 8'sd66}, {11'sd897, 10'sd505, 11'sd593}, {11'sd918, 9'sd232, 11'sd-926}},
{{13'sd-2293, 12'sd1152, 12'sd1488}, {13'sd2502, 10'sd441, 12'sd-1664}, {12'sd1083, 10'sd354, 13'sd-2063}},
{{13'sd-2764, 12'sd1411, 12'sd-1440}, {12'sd-1154, 12'sd1723, 11'sd-696}, {13'sd-2240, 12'sd-1365, 12'sd-1709}},
{{12'sd1653, 9'sd196, 12'sd-1819}, {9'sd-168, 12'sd1217, 12'sd-1767}, {13'sd-2098, 13'sd-2196, 12'sd-1638}},
{{11'sd-586, 13'sd2622, 13'sd2188}, {11'sd-601, 9'sd185, 11'sd924}, {11'sd932, 10'sd-469, 12'sd-2036}},
{{12'sd-2018, 12'sd-1416, 11'sd890}, {12'sd1812, 11'sd998, 13'sd-3510}, {13'sd-2856, 12'sd1498, 11'sd907}},
{{12'sd1828, 9'sd-133, 11'sd514}, {12'sd1431, 12'sd-1960, 8'sd-107}, {11'sd-744, 12'sd1205, 9'sd187}},
{{12'sd-1858, 7'sd-61, 9'sd129}, {13'sd2382, 13'sd-2464, 10'sd-408}, {10'sd-375, 12'sd-1684, 13'sd2322}},
{{13'sd-2433, 6'sd-31, 12'sd-1344}, {8'sd94, 10'sd458, 11'sd-621}, {12'sd-1224, 11'sd729, 13'sd-2075}},
{{8'sd-64, 13'sd2616, 12'sd-1234}, {9'sd189, 12'sd2033, 11'sd-546}, {9'sd-241, 12'sd-1524, 12'sd1535}},
{{9'sd-141, 7'sd53, 10'sd400}, {12'sd-1168, 13'sd2163, 13'sd2237}, {12'sd1903, 12'sd-1834, 12'sd-1797}},
{{10'sd278, 13'sd-2546, 12'sd1040}, {13'sd2146, 11'sd809, 13'sd2595}, {9'sd255, 13'sd2691, 12'sd1640}},
{{12'sd2013, 12'sd1253, 12'sd-1982}, {13'sd2154, 10'sd-499, 13'sd-2156}, {12'sd-1033, 11'sd-579, 10'sd-258}},
{{13'sd2750, 12'sd-1056, 13'sd2597}, {13'sd2161, 11'sd-876, 10'sd-508}, {10'sd342, 13'sd-2415, 13'sd-2118}},
{{13'sd2630, 10'sd-358, 12'sd-1322}, {6'sd16, 12'sd-1502, 13'sd2729}, {13'sd-2227, 11'sd688, 12'sd1183}},
{{13'sd-2229, 13'sd-2456, 8'sd93}, {11'sd952, 12'sd-1468, 10'sd-463}, {13'sd-2420, 10'sd-452, 12'sd1913}},
{{9'sd-223, 11'sd815, 11'sd622}, {8'sd119, 12'sd1929, 9'sd-228}, {12'sd1883, 12'sd-1518, 11'sd-839}},
{{11'sd768, 12'sd1811, 12'sd1360}, {13'sd2822, 12'sd1966, 10'sd460}, {13'sd2129, 12'sd-1409, 7'sd-36}},
{{12'sd-2006, 11'sd908, 11'sd1019}, {7'sd51, 11'sd736, 13'sd-2072}, {11'sd-648, 11'sd-908, 12'sd1683}},
{{12'sd1721, 10'sd449, 11'sd545}, {12'sd1046, 13'sd2424, 12'sd-1749}, {12'sd-1974, 8'sd-110, 13'sd2933}},
{{10'sd347, 10'sd289, 9'sd216}, {11'sd645, 13'sd2346, 9'sd201}, {9'sd230, 12'sd-1146, 10'sd329}},
{{10'sd-490, 11'sd870, 12'sd-2037}, {12'sd-1855, 12'sd-1630, 12'sd-1437}, {12'sd-1137, 11'sd-1020, 12'sd-1355}},
{{9'sd218, 13'sd2090, 12'sd-1132}, {11'sd-909, 7'sd-50, 11'sd520}, {11'sd913, 13'sd2420, 12'sd1294}},
{{13'sd-2334, 12'sd1935, 10'sd-407}, {12'sd1311, 11'sd712, 11'sd-646}, {13'sd-2222, 12'sd1215, 12'sd1923}},
{{12'sd1710, 12'sd-1097, 13'sd3119}, {12'sd1797, 12'sd1647, 10'sd272}, {11'sd591, 11'sd-910, 12'sd1150}},
{{13'sd-2523, 13'sd-2811, 12'sd1183}, {12'sd-1976, 11'sd-778, 13'sd-2205}, {13'sd-2896, 12'sd1583, 12'sd1296}},
{{12'sd-1421, 12'sd-1486, 12'sd-1127}, {13'sd2523, 12'sd1480, 11'sd668}, {12'sd-1886, 13'sd2706, 11'sd-569}},
{{11'sd583, 13'sd-2519, 7'sd-50}, {12'sd-1994, 13'sd2506, 13'sd2641}, {11'sd-1000, 11'sd988, 12'sd1465}},
{{13'sd-2104, 12'sd-1411, 13'sd-2102}, {11'sd-675, 11'sd-711, 12'sd-1889}, {13'sd-2160, 11'sd-531, 13'sd-3655}},
{{9'sd-217, 12'sd1809, 11'sd-643}, {12'sd1513, 11'sd-714, 12'sd1206}, {6'sd30, 13'sd2104, 12'sd-1242}},
{{12'sd-1460, 12'sd1545, 13'sd-2088}, {12'sd1555, 10'sd300, 12'sd1146}, {13'sd2277, 12'sd1307, 13'sd3011}},
{{13'sd3205, 13'sd2128, 13'sd2084}, {11'sd541, 8'sd125, 13'sd-2109}, {12'sd-1757, 10'sd470, 10'sd319}},
{{10'sd-392, 13'sd-2260, 12'sd-1979}, {10'sd-269, 11'sd-693, 12'sd-1114}, {13'sd2135, 13'sd2599, 12'sd2033}},
{{10'sd-493, 13'sd2158, 13'sd2173}, {12'sd1058, 13'sd-2054, 6'sd19}, {12'sd1867, 13'sd2323, 10'sd-258}},
{{12'sd-1584, 12'sd1455, 12'sd1294}, {5'sd-11, 12'sd1763, 11'sd-620}, {12'sd-1567, 13'sd-2488, 13'sd2668}},
{{10'sd317, 13'sd-2178, 12'sd-1325}, {11'sd715, 11'sd-648, 12'sd1096}, {13'sd-2221, 10'sd-503, 12'sd1832}},
{{10'sd-402, 12'sd2031, 8'sd109}, {11'sd-938, 13'sd2211, 12'sd1126}, {12'sd1502, 12'sd-1806, 10'sd-479}},
{{11'sd-598, 12'sd1315, 13'sd2215}, {12'sd1107, 12'sd1893, 12'sd-1310}, {12'sd-1903, 11'sd-795, 11'sd931}},
{{9'sd251, 12'sd1730, 12'sd1881}, {13'sd-2611, 12'sd-1833, 12'sd-1096}, {11'sd-625, 10'sd302, 12'sd-1881}},
{{13'sd-2084, 10'sd-326, 12'sd-1551}, {12'sd1127, 13'sd2661, 11'sd-663}, {10'sd418, 11'sd-717, 12'sd-1886}},
{{13'sd-2506, 10'sd277, 11'sd733}, {12'sd-1377, 12'sd1311, 12'sd-1027}, {13'sd2920, 10'sd-369, 12'sd-1466}},
{{12'sd1562, 9'sd213, 12'sd1584}, {13'sd2392, 12'sd-2045, 12'sd-1430}, {9'sd251, 12'sd1292, 13'sd-2325}},
{{11'sd838, 11'sd970, 9'sd-226}, {12'sd1901, 12'sd-1611, 12'sd1573}, {13'sd-2362, 12'sd-1245, 9'sd-139}},
{{12'sd1727, 12'sd-1045, 11'sd771}, {2'sd1, 13'sd2246, 12'sd1279}, {10'sd303, 12'sd1677, 13'sd2065}},
{{13'sd-3448, 10'sd-398, 13'sd-3414}, {11'sd-661, 12'sd-2018, 9'sd-231}, {12'sd1628, 13'sd2604, 11'sd-829}},
{{11'sd905, 4'sd-4, 12'sd1883}, {13'sd-2592, 10'sd436, 11'sd963}, {12'sd-1401, 13'sd-2589, 13'sd-3114}},
{{13'sd2626, 13'sd2131, 11'sd684}, {11'sd-856, 12'sd1943, 13'sd-2183}, {9'sd-129, 12'sd1434, 12'sd-1630}},
{{11'sd739, 10'sd404, 10'sd474}, {12'sd1149, 11'sd528, 12'sd1113}, {12'sd-1836, 6'sd-22, 11'sd1006}},
{{12'sd-1438, 12'sd1769, 12'sd-1612}, {12'sd-1260, 11'sd607, 11'sd-993}, {12'sd1355, 13'sd-2527, 13'sd-3020}},
{{12'sd-1780, 13'sd-2616, 13'sd-2255}, {12'sd-1177, 12'sd-1695, 11'sd928}, {12'sd1517, 12'sd-1773, 12'sd1696}},
{{11'sd683, 12'sd-1520, 13'sd2100}, {11'sd677, 9'sd129, 9'sd-172}, {11'sd-961, 12'sd-1333, 11'sd-531}},
{{13'sd3368, 13'sd2125, 11'sd915}, {13'sd2071, 12'sd1041, 11'sd579}, {13'sd2444, 12'sd1393, 11'sd-891}}},
{
{{8'sd-106, 12'sd1939, 12'sd-1826}, {10'sd274, 11'sd853, 11'sd550}, {12'sd-1726, 13'sd2081, 12'sd-1696}},
{{11'sd-766, 12'sd-1207, 13'sd-2281}, {10'sd-281, 12'sd1343, 12'sd1549}, {12'sd1703, 12'sd-1416, 8'sd100}},
{{13'sd2393, 11'sd1011, 12'sd1185}, {11'sd721, 11'sd-685, 12'sd1698}, {12'sd1848, 13'sd-2110, 9'sd236}},
{{7'sd-39, 8'sd-81, 9'sd200}, {11'sd-851, 9'sd-213, 11'sd-842}, {13'sd2432, 11'sd-805, 11'sd634}},
{{10'sd-417, 10'sd-344, 10'sd-256}, {12'sd1220, 4'sd6, 12'sd1106}, {12'sd1549, 11'sd654, 10'sd431}},
{{11'sd-623, 13'sd-2913, 11'sd581}, {12'sd1434, 11'sd-1020, 9'sd247}, {12'sd-1795, 12'sd1347, 12'sd2034}},
{{13'sd2676, 11'sd-975, 13'sd2048}, {12'sd1209, 9'sd200, 8'sd71}, {13'sd2186, 11'sd-888, 12'sd1175}},
{{12'sd1451, 13'sd2404, 12'sd1983}, {11'sd-654, 13'sd2882, 9'sd-169}, {10'sd270, 11'sd850, 13'sd-2112}},
{{9'sd-138, 12'sd1430, 13'sd-2238}, {12'sd-1380, 13'sd-2204, 12'sd-1447}, {11'sd-657, 13'sd2548, 11'sd-602}},
{{12'sd1189, 13'sd2277, 12'sd-1154}, {13'sd-2573, 12'sd1876, 13'sd3041}, {12'sd-1141, 13'sd3193, 13'sd2397}},
{{13'sd2376, 12'sd1419, 12'sd1857}, {11'sd-534, 10'sd309, 12'sd-1308}, {10'sd467, 12'sd-1130, 12'sd-1033}},
{{13'sd2431, 12'sd-1804, 6'sd28}, {12'sd1246, 12'sd-1118, 13'sd-2994}, {13'sd-2273, 11'sd-775, 12'sd1127}},
{{12'sd-1372, 11'sd-662, 12'sd-1101}, {11'sd-720, 11'sd970, 12'sd-1532}, {10'sd305, 11'sd-1007, 11'sd566}},
{{12'sd-1385, 11'sd652, 11'sd-850}, {12'sd-1050, 13'sd-2168, 12'sd-1224}, {11'sd-777, 9'sd-217, 12'sd-1676}},
{{8'sd-93, 13'sd-2229, 12'sd1448}, {11'sd850, 11'sd-526, 13'sd2614}, {13'sd2575, 13'sd2718, 12'sd1106}},
{{8'sd-93, 12'sd-1430, 12'sd-1929}, {11'sd929, 12'sd-1981, 12'sd1847}, {12'sd-1624, 8'sd95, 10'sd308}},
{{12'sd1424, 12'sd-1464, 13'sd-2183}, {13'sd2296, 13'sd-2615, 12'sd1067}, {12'sd-1929, 12'sd-2036, 11'sd-1014}},
{{13'sd2607, 11'sd618, 13'sd2702}, {7'sd-54, 11'sd820, 13'sd2088}, {12'sd-1064, 12'sd1866, 10'sd-276}},
{{12'sd-1914, 12'sd1159, 13'sd2108}, {12'sd1473, 12'sd2030, 10'sd-424}, {12'sd1647, 12'sd-1841, 12'sd1532}},
{{11'sd570, 8'sd-119, 13'sd2668}, {13'sd-2789, 12'sd2000, 11'sd-903}, {11'sd-593, 10'sd-457, 12'sd-1269}},
{{13'sd2098, 13'sd-2508, 12'sd1202}, {12'sd-1853, 12'sd1464, 12'sd-1577}, {12'sd1612, 12'sd-1583, 12'sd-1382}},
{{12'sd1857, 12'sd-1250, 12'sd1625}, {10'sd361, 12'sd1311, 12'sd-1369}, {12'sd-1969, 12'sd1664, 11'sd-989}},
{{12'sd-1113, 10'sd-299, 12'sd1307}, {11'sd542, 13'sd2744, 12'sd1307}, {13'sd2362, 13'sd2869, 11'sd659}},
{{12'sd-1650, 12'sd-1038, 12'sd1241}, {12'sd1480, 12'sd-1981, 13'sd2994}, {11'sd568, 13'sd2349, 11'sd-847}},
{{11'sd536, 13'sd-2317, 12'sd1242}, {13'sd2322, 7'sd33, 13'sd2362}, {9'sd207, 12'sd-1145, 11'sd-631}},
{{13'sd2678, 10'sd-411, 12'sd1838}, {12'sd1246, 10'sd260, 11'sd607}, {12'sd1813, 12'sd-1129, 10'sd291}},
{{10'sd-316, 13'sd-2242, 11'sd-787}, {10'sd-395, 13'sd-2351, 12'sd1235}, {12'sd1787, 11'sd-688, 10'sd-474}},
{{13'sd-2820, 13'sd-2943, 10'sd351}, {13'sd2130, 12'sd-1630, 12'sd-1241}, {12'sd1157, 9'sd238, 12'sd-1199}},
{{13'sd-2190, 11'sd-669, 11'sd-993}, {12'sd1159, 12'sd2041, 7'sd-45}, {12'sd1143, 12'sd-1906, 13'sd2642}},
{{11'sd-1023, 12'sd1893, 9'sd-162}, {13'sd2074, 11'sd-609, 12'sd1345}, {10'sd-441, 11'sd-948, 13'sd-2979}},
{{10'sd260, 9'sd-130, 13'sd2428}, {13'sd-2235, 12'sd1854, 10'sd410}, {12'sd-1636, 9'sd176, 11'sd-834}},
{{12'sd-1848, 12'sd1322, 12'sd-1599}, {12'sd1314, 13'sd2261, 13'sd2638}, {13'sd-2826, 12'sd-1584, 12'sd1810}},
{{13'sd-2591, 12'sd1077, 11'sd-530}, {12'sd-1543, 12'sd1721, 9'sd-216}, {12'sd-2047, 12'sd1175, 13'sd2448}},
{{12'sd-1638, 9'sd237, 12'sd1332}, {11'sd-519, 12'sd1940, 10'sd377}, {13'sd-2187, 12'sd1804, 13'sd-2375}},
{{12'sd1582, 13'sd-2192, 12'sd1318}, {12'sd1450, 8'sd-110, 8'sd118}, {12'sd1661, 9'sd-156, 11'sd-735}},
{{11'sd-966, 13'sd2342, 11'sd706}, {12'sd1434, 10'sd393, 13'sd2368}, {13'sd2140, 13'sd2054, 11'sd-894}},
{{12'sd-1940, 12'sd-1411, 13'sd-2913}, {9'sd185, 13'sd-2940, 7'sd45}, {10'sd261, 11'sd710, 12'sd1535}},
{{11'sd609, 12'sd-1652, 12'sd1767}, {10'sd-310, 11'sd-839, 12'sd1311}, {12'sd-1055, 6'sd-26, 10'sd290}},
{{13'sd-2359, 11'sd687, 11'sd600}, {13'sd-2140, 12'sd1960, 11'sd971}, {13'sd2574, 10'sd-285, 12'sd1852}},
{{12'sd1380, 11'sd1016, 11'sd-740}, {11'sd821, 12'sd-1776, 12'sd1828}, {12'sd1492, 13'sd-2513, 11'sd742}},
{{12'sd-2005, 12'sd1688, 11'sd-900}, {13'sd-2307, 4'sd5, 12'sd1182}, {13'sd2229, 12'sd1970, 11'sd536}},
{{13'sd-2251, 13'sd-2379, 12'sd1141}, {9'sd171, 12'sd-1175, 12'sd1186}, {11'sd699, 6'sd28, 12'sd1175}},
{{13'sd2068, 13'sd-2226, 11'sd594}, {11'sd-955, 13'sd2999, 13'sd-2158}, {10'sd284, 12'sd-1522, 8'sd125}},
{{13'sd-3362, 13'sd-2091, 11'sd-825}, {13'sd2110, 13'sd-2471, 13'sd-3284}, {14'sd-4584, 9'sd142, 10'sd370}},
{{12'sd-1529, 12'sd1572, 9'sd-154}, {12'sd-1777, 9'sd193, 12'sd1706}, {10'sd-274, 12'sd-1660, 11'sd-641}},
{{12'sd2046, 12'sd-1587, 11'sd-541}, {12'sd-1617, 12'sd-1474, 13'sd-2450}, {12'sd-1293, 13'sd-2066, 9'sd-160}},
{{10'sd-395, 12'sd1503, 13'sd-2415}, {12'sd-1751, 11'sd888, 12'sd-1686}, {9'sd237, 9'sd-216, 13'sd-2427}},
{{13'sd2204, 12'sd1909, 12'sd1067}, {11'sd616, 10'sd-510, 12'sd1776}, {13'sd2153, 12'sd-1831, 12'sd1482}},
{{13'sd2432, 12'sd1797, 13'sd-3678}, {12'sd-1957, 12'sd1184, 10'sd-458}, {12'sd1993, 12'sd1326, 11'sd933}},
{{13'sd2935, 12'sd1100, 13'sd-2326}, {13'sd-2375, 11'sd856, 13'sd-2181}, {13'sd2241, 12'sd-1733, 13'sd-2089}},
{{12'sd1312, 9'sd190, 12'sd-1949}, {12'sd-1474, 7'sd49, 12'sd-1403}, {12'sd-1358, 8'sd-78, 11'sd542}},
{{12'sd2031, 12'sd1172, 13'sd2262}, {10'sd-452, 9'sd-139, 11'sd533}, {11'sd-1018, 10'sd-405, 12'sd1839}},
{{12'sd-1090, 13'sd2357, 12'sd1415}, {12'sd-1538, 10'sd-457, 9'sd147}, {13'sd-2388, 12'sd1851, 11'sd-908}},
{{12'sd1480, 13'sd2910, 11'sd-933}, {12'sd1049, 11'sd-628, 12'sd-1932}, {12'sd-1377, 11'sd-818, 13'sd2720}},
{{13'sd2553, 13'sd2785, 10'sd-296}, {12'sd-1066, 12'sd-1279, 13'sd-2087}, {11'sd866, 11'sd753, 13'sd2690}},
{{12'sd-1083, 9'sd-192, 12'sd-1971}, {11'sd568, 9'sd-137, 12'sd-1531}, {13'sd2616, 9'sd-205, 13'sd2332}},
{{9'sd222, 12'sd-1317, 13'sd2053}, {13'sd2250, 12'sd-1131, 13'sd2270}, {13'sd2670, 13'sd3226, 12'sd2003}},
{{9'sd-146, 11'sd900, 10'sd316}, {10'sd-404, 12'sd1974, 12'sd1538}, {13'sd2639, 12'sd-1863, 12'sd-1721}},
{{12'sd1826, 10'sd-409, 12'sd1450}, {12'sd1419, 13'sd-2202, 11'sd740}, {12'sd-1597, 12'sd-1478, 13'sd2486}},
{{13'sd3507, 12'sd1973, 12'sd1790}, {12'sd2044, 12'sd-1712, 13'sd2305}, {11'sd782, 11'sd783, 10'sd330}},
{{10'sd358, 11'sd-691, 13'sd-2153}, {12'sd-1851, 11'sd-615, 13'sd2230}, {6'sd-25, 12'sd-1906, 12'sd1574}},
{{11'sd824, 11'sd-812, 13'sd-2369}, {12'sd1408, 12'sd-1194, 10'sd-384}, {13'sd2835, 13'sd-2639, 10'sd-500}},
{{12'sd1078, 12'sd-1066, 11'sd595}, {11'sd810, 10'sd-323, 13'sd-2391}, {9'sd-163, 13'sd2461, 13'sd2363}},
{{13'sd-3366, 12'sd1443, 10'sd-409}, {13'sd-2318, 12'sd-1822, 12'sd-1305}, {11'sd-752, 12'sd1776, 12'sd-1933}}},
{
{{13'sd2638, 12'sd-1754, 13'sd-2683}, {12'sd1642, 12'sd1626, 12'sd-1793}, {13'sd2193, 10'sd478, 12'sd-1114}},
{{12'sd1069, 13'sd-2623, 13'sd2084}, {12'sd1235, 11'sd617, 11'sd-678}, {11'sd-639, 13'sd2215, 12'sd-1619}},
{{12'sd1361, 11'sd-650, 12'sd1838}, {12'sd1789, 10'sd-422, 13'sd2311}, {11'sd-729, 13'sd2287, 12'sd-1621}},
{{12'sd-1314, 12'sd1772, 12'sd1717}, {12'sd1591, 12'sd1863, 13'sd-2853}, {12'sd-2017, 13'sd-2524, 10'sd300}},
{{13'sd3485, 13'sd2870, 6'sd16}, {11'sd624, 12'sd1106, 13'sd-3623}, {12'sd-1504, 12'sd1231, 13'sd-3909}},
{{11'sd-552, 12'sd1849, 11'sd-546}, {13'sd2672, 12'sd-1363, 13'sd-3625}, {10'sd-462, 11'sd533, 13'sd-2424}},
{{13'sd-2240, 12'sd1819, 14'sd-4629}, {12'sd1446, 11'sd-548, 13'sd-3871}, {12'sd-1317, 12'sd-1601, 11'sd634}},
{{11'sd-625, 11'sd549, 13'sd-2856}, {12'sd-1536, 9'sd135, 10'sd-508}, {12'sd1424, 12'sd1579, 8'sd112}},
{{12'sd1497, 9'sd247, 13'sd-2160}, {10'sd458, 12'sd-1797, 10'sd-331}, {12'sd1851, 12'sd1340, 13'sd-2639}},
{{12'sd-1128, 11'sd-686, 9'sd-217}, {12'sd1868, 10'sd-442, 11'sd1010}, {13'sd2685, 13'sd2656, 13'sd-2426}},
{{12'sd-1061, 10'sd-256, 13'sd2538}, {12'sd-1181, 12'sd1141, 13'sd-2708}, {12'sd1097, 13'sd2563, 8'sd-68}},
{{11'sd1018, 12'sd-1319, 13'sd2215}, {12'sd1490, 13'sd2736, 13'sd2137}, {13'sd-2765, 10'sd-303, 13'sd-2739}},
{{13'sd2119, 10'sd319, 11'sd536}, {12'sd1837, 12'sd-1627, 11'sd746}, {12'sd-1156, 11'sd-776, 8'sd-83}},
{{11'sd811, 13'sd-2497, 9'sd172}, {7'sd46, 9'sd233, 11'sd-992}, {12'sd-2030, 12'sd1503, 13'sd2050}},
{{11'sd596, 12'sd1093, 13'sd-2208}, {11'sd853, 11'sd650, 13'sd-2386}, {11'sd-997, 10'sd257, 11'sd-908}},
{{13'sd2230, 12'sd-1231, 9'sd186}, {13'sd-2360, 13'sd-2390, 11'sd1016}, {12'sd-1588, 11'sd662, 11'sd787}},
{{13'sd-2339, 13'sd-2877, 12'sd1589}, {10'sd-428, 12'sd1238, 11'sd788}, {10'sd468, 11'sd-589, 11'sd753}},
{{12'sd1915, 13'sd-2224, 13'sd-2214}, {12'sd1977, 11'sd598, 12'sd1125}, {13'sd-2668, 11'sd645, 11'sd844}},
{{12'sd-1163, 10'sd489, 10'sd422}, {12'sd-1971, 12'sd1614, 12'sd-2017}, {10'sd437, 13'sd-2240, 13'sd2788}},
{{12'sd1695, 12'sd1184, 13'sd-2108}, {12'sd-1623, 12'sd1636, 13'sd3400}, {11'sd-956, 12'sd-1298, 12'sd-1095}},
{{12'sd-1242, 13'sd-2770, 8'sd76}, {13'sd-2793, 13'sd-2696, 9'sd146}, {11'sd-898, 13'sd-2239, 13'sd-2270}},
{{13'sd-2594, 12'sd1446, 12'sd1301}, {12'sd1712, 9'sd233, 13'sd2832}, {10'sd385, 12'sd1550, 11'sd696}},
{{12'sd1344, 12'sd-1881, 10'sd364}, {12'sd-1914, 7'sd-57, 12'sd1561}, {12'sd-1284, 12'sd1551, 11'sd-561}},
{{10'sd-444, 12'sd1633, 12'sd-1121}, {11'sd-740, 12'sd1705, 12'sd2039}, {12'sd-1806, 10'sd-359, 13'sd3527}},
{{10'sd-465, 9'sd-252, 5'sd-11}, {13'sd2470, 12'sd-1433, 12'sd1925}, {12'sd-1902, 10'sd-471, 13'sd2253}},
{{11'sd-944, 12'sd1907, 12'sd-1138}, {10'sd473, 12'sd-1595, 10'sd501}, {12'sd-1309, 9'sd-166, 13'sd-2730}},
{{11'sd-741, 10'sd-355, 13'sd2199}, {10'sd-270, 10'sd-330, 10'sd440}, {11'sd-592, 11'sd639, 12'sd-1402}},
{{13'sd2670, 8'sd105, 13'sd-2306}, {13'sd-2745, 13'sd-2477, 12'sd-1545}, {12'sd-1540, 9'sd-135, 12'sd1039}},
{{13'sd3084, 12'sd-1593, 9'sd-206}, {12'sd-1698, 12'sd-1321, 9'sd212}, {12'sd1700, 8'sd-123, 13'sd3938}},
{{11'sd778, 12'sd-1561, 13'sd2298}, {13'sd2334, 12'sd1195, 13'sd2596}, {13'sd3073, 12'sd-1411, 9'sd-190}},
{{12'sd-1080, 12'sd-1319, 12'sd-1365}, {13'sd-2161, 11'sd-586, 13'sd2807}, {12'sd-1038, 13'sd-2395, 13'sd2594}},
{{12'sd1614, 13'sd3353, 12'sd1419}, {11'sd-516, 10'sd-379, 12'sd-1681}, {9'sd140, 10'sd-273, 13'sd-2320}},
{{11'sd-822, 11'sd715, 12'sd-1774}, {12'sd-1615, 10'sd-328, 10'sd418}, {9'sd178, 12'sd-1071, 11'sd941}},
{{13'sd3705, 11'sd595, 12'sd-1419}, {13'sd2358, 12'sd-1423, 12'sd-1248}, {11'sd-994, 9'sd128, 11'sd759}},
{{12'sd-1364, 11'sd-915, 10'sd-461}, {12'sd1064, 11'sd547, 11'sd928}, {13'sd-2739, 10'sd458, 12'sd-1176}},
{{11'sd-758, 12'sd-1129, 10'sd267}, {13'sd2375, 11'sd664, 9'sd-229}, {13'sd2281, 12'sd-1462, 12'sd-1329}},
{{13'sd-3164, 11'sd-990, 12'sd-1060}, {12'sd-1376, 2'sd1, 10'sd-347}, {14'sd-5390, 13'sd-2794, 11'sd937}},
{{13'sd2980, 13'sd-2939, 13'sd2067}, {13'sd-2491, 11'sd519, 11'sd543}, {7'sd-48, 12'sd1111, 13'sd-2614}},
{{12'sd1909, 10'sd-477, 13'sd2309}, {13'sd-2454, 12'sd-1995, 12'sd-1754}, {12'sd1164, 12'sd1556, 13'sd-2146}},
{{12'sd-1679, 12'sd-1179, 13'sd-2105}, {12'sd-1502, 11'sd827, 13'sd-2691}, {11'sd-669, 13'sd2167, 13'sd-2499}},
{{12'sd-1631, 12'sd-1614, 12'sd1086}, {12'sd-1242, 12'sd1106, 13'sd-2629}, {10'sd-261, 12'sd-1854, 12'sd-2029}},
{{12'sd1224, 11'sd-557, 12'sd-1949}, {11'sd1008, 13'sd-2583, 13'sd-2500}, {12'sd1526, 10'sd-458, 13'sd-2654}},
{{12'sd1555, 11'sd875, 13'sd-2853}, {9'sd-199, 13'sd2528, 9'sd-128}, {12'sd-1024, 12'sd1778, 6'sd23}},
{{13'sd2260, 10'sd453, 11'sd-897}, {13'sd2056, 13'sd-2738, 12'sd-1996}, {7'sd-36, 11'sd695, 13'sd-3329}},
{{12'sd-1940, 12'sd1288, 13'sd-2485}, {13'sd-2148, 10'sd-361, 9'sd252}, {13'sd2455, 11'sd795, 8'sd-98}},
{{13'sd-2614, 11'sd955, 12'sd-1092}, {13'sd2130, 13'sd-2178, 9'sd-193}, {11'sd-586, 6'sd24, 12'sd1411}},
{{13'sd-2087, 10'sd-320, 12'sd-1101}, {12'sd-1162, 13'sd2098, 12'sd2006}, {13'sd-2744, 12'sd2027, 13'sd2612}},
{{10'sd-383, 12'sd1624, 12'sd1793}, {11'sd627, 11'sd-642, 13'sd2243}, {10'sd345, 11'sd757, 13'sd2663}},
{{13'sd2265, 12'sd1451, 11'sd-982}, {12'sd1849, 12'sd1892, 11'sd684}, {11'sd669, 11'sd556, 9'sd197}},
{{14'sd-4541, 13'sd-3362, 8'sd-108}, {12'sd-1835, 13'sd2092, 11'sd-961}, {13'sd-3656, 6'sd-27, 13'sd2380}},
{{13'sd3112, 8'sd92, 13'sd2091}, {11'sd667, 12'sd1290, 13'sd2091}, {12'sd-1844, 12'sd1382, 12'sd1742}},
{{12'sd-1373, 13'sd2600, 12'sd-1149}, {8'sd76, 13'sd2196, 11'sd1021}, {11'sd-906, 13'sd-2232, 12'sd-1424}},
{{7'sd60, 12'sd-1826, 11'sd-654}, {12'sd-1454, 11'sd999, 10'sd385}, {12'sd2029, 13'sd3377, 12'sd-1125}},
{{10'sd303, 9'sd-140, 13'sd2337}, {12'sd1547, 11'sd640, 13'sd2486}, {13'sd-2316, 11'sd696, 11'sd594}},
{{11'sd762, 11'sd871, 13'sd-3130}, {12'sd-1786, 12'sd-1325, 11'sd724}, {9'sd-139, 11'sd745, 14'sd-4968}},
{{11'sd-1013, 12'sd1445, 13'sd-2270}, {12'sd-1221, 13'sd-2486, 12'sd-1544}, {11'sd-884, 13'sd-2537, 11'sd889}},
{{11'sd850, 13'sd-2912, 13'sd-2717}, {6'sd17, 10'sd-444, 14'sd-4359}, {12'sd-1298, 13'sd-2510, 11'sd570}},
{{11'sd-796, 12'sd1710, 12'sd1662}, {11'sd-650, 12'sd-1046, 13'sd-2293}, {8'sd-66, 11'sd949, 12'sd-2043}},
{{12'sd1845, 9'sd-218, 13'sd-3125}, {10'sd302, 12'sd-1737, 12'sd1636}, {10'sd267, 13'sd-2137, 10'sd-486}},
{{12'sd1085, 13'sd3760, 11'sd630}, {12'sd-1521, 13'sd3500, 11'sd986}, {11'sd565, 11'sd851, 7'sd-60}},
{{12'sd1911, 11'sd655, 13'sd2574}, {10'sd-346, 12'sd-1586, 13'sd2775}, {12'sd-1963, 13'sd-2940, 8'sd121}},
{{13'sd2726, 9'sd-171, 11'sd-519}, {13'sd2158, 11'sd-957, 13'sd-2577}, {11'sd-639, 9'sd245, 13'sd-3834}},
{{14'sd-4125, 12'sd1086, 13'sd-2153}, {13'sd-2835, 13'sd-3994, 10'sd-407}, {11'sd-866, 13'sd-3066, 11'sd973}},
{{12'sd1319, 12'sd1216, 12'sd-1862}, {9'sd133, 12'sd1547, 11'sd968}, {13'sd3388, 12'sd1431, 12'sd1049}}},
{
{{12'sd-1128, 8'sd-108, 12'sd-1188}, {12'sd-1766, 12'sd-1531, 12'sd1027}, {12'sd-1110, 10'sd-292, 12'sd1890}},
{{13'sd-2638, 11'sd-730, 11'sd-856}, {13'sd2636, 12'sd1552, 12'sd1484}, {12'sd-1400, 12'sd1861, 12'sd1762}},
{{12'sd1968, 12'sd-1882, 12'sd1674}, {13'sd2225, 11'sd675, 13'sd2065}, {9'sd150, 12'sd1318, 12'sd1545}},
{{12'sd1066, 11'sd727, 12'sd-1567}, {12'sd1686, 12'sd-1104, 12'sd1985}, {12'sd1329, 12'sd1749, 10'sd409}},
{{12'sd1712, 13'sd2340, 12'sd1236}, {11'sd-752, 12'sd-1555, 11'sd608}, {13'sd-3088, 13'sd-2246, 9'sd169}},
{{13'sd2475, 11'sd681, 9'sd249}, {13'sd-2203, 12'sd1103, 9'sd-196}, {10'sd405, 12'sd1423, 12'sd1425}},
{{11'sd-969, 11'sd956, 11'sd-693}, {11'sd-760, 9'sd174, 12'sd1029}, {11'sd688, 13'sd-2703, 10'sd329}},
{{11'sd-895, 11'sd519, 12'sd1337}, {10'sd455, 9'sd169, 13'sd2438}, {9'sd-194, 11'sd-956, 13'sd2601}},
{{13'sd2106, 12'sd-1813, 9'sd199}, {12'sd1860, 11'sd-944, 12'sd-1779}, {13'sd-2051, 12'sd-1728, 12'sd1154}},
{{12'sd-1097, 10'sd-397, 12'sd1409}, {13'sd2279, 12'sd-1564, 11'sd916}, {13'sd-2123, 10'sd319, 10'sd361}},
{{9'sd-231, 12'sd-1663, 10'sd-444}, {11'sd-683, 6'sd-31, 13'sd-2391}, {13'sd2606, 12'sd-1596, 12'sd1211}},
{{12'sd1549, 12'sd1469, 12'sd1873}, {12'sd1252, 11'sd905, 11'sd975}, {10'sd316, 11'sd743, 11'sd-862}},
{{10'sd364, 12'sd1861, 12'sd1826}, {13'sd2889, 12'sd-1973, 12'sd-2003}, {11'sd749, 10'sd469, 12'sd1595}},
{{13'sd2051, 11'sd598, 9'sd-245}, {13'sd-2738, 10'sd-258, 11'sd-680}, {12'sd-1519, 11'sd753, 11'sd729}},
{{13'sd-2681, 11'sd-593, 13'sd-3409}, {13'sd2462, 12'sd-1967, 11'sd627}, {12'sd-1464, 12'sd-2017, 13'sd-2573}},
{{12'sd1585, 12'sd1706, 13'sd2069}, {13'sd2511, 12'sd1268, 11'sd519}, {12'sd1186, 11'sd533, 13'sd2322}},
{{12'sd-1757, 13'sd2511, 9'sd131}, {12'sd-1579, 12'sd1245, 11'sd-824}, {9'sd-173, 10'sd413, 11'sd612}},
{{11'sd816, 12'sd-1737, 12'sd-1342}, {11'sd-774, 13'sd-2109, 12'sd1789}, {11'sd977, 13'sd2396, 13'sd2712}},
{{11'sd529, 10'sd377, 11'sd-824}, {9'sd243, 12'sd1133, 12'sd-1357}, {13'sd2184, 9'sd-207, 13'sd-2053}},
{{10'sd-310, 12'sd1038, 13'sd2095}, {13'sd-2108, 12'sd-1581, 13'sd-2594}, {12'sd1923, 12'sd-1179, 12'sd-1548}},
{{13'sd-2366, 13'sd2261, 13'sd-2745}, {12'sd-1341, 12'sd1104, 11'sd-1008}, {6'sd23, 13'sd-2229, 9'sd152}},
{{9'sd-207, 12'sd-1472, 11'sd-1002}, {12'sd1729, 12'sd-1860, 12'sd1446}, {12'sd1114, 13'sd-2714, 13'sd2439}},
{{12'sd-1666, 11'sd-594, 10'sd386}, {11'sd-578, 13'sd-2630, 10'sd-407}, {12'sd-1111, 10'sd271, 11'sd-532}},
{{13'sd-2542, 11'sd-670, 13'sd2768}, {8'sd97, 13'sd-2248, 13'sd2805}, {13'sd2533, 12'sd1100, 9'sd201}},
{{11'sd926, 12'sd1140, 10'sd-307}, {11'sd-910, 8'sd108, 12'sd-1649}, {10'sd362, 12'sd-1377, 12'sd1122}},
{{13'sd2335, 12'sd-1422, 12'sd-1964}, {11'sd-796, 12'sd-1243, 12'sd-1323}, {12'sd1884, 12'sd-1973, 10'sd268}},
{{13'sd2435, 13'sd2856, 9'sd-158}, {11'sd-908, 8'sd-78, 11'sd970}, {14'sd4230, 9'sd-148, 8'sd79}},
{{13'sd-2223, 10'sd-296, 13'sd-2688}, {13'sd2593, 8'sd-93, 12'sd1024}, {9'sd133, 12'sd1284, 12'sd-1621}},
{{10'sd-431, 10'sd-404, 13'sd-2350}, {10'sd352, 10'sd-410, 9'sd170}, {7'sd-38, 13'sd2494, 11'sd-665}},
{{12'sd1926, 11'sd-805, 11'sd-1012}, {12'sd-1115, 13'sd3079, 12'sd1868}, {10'sd372, 12'sd-1123, 9'sd-129}},
{{9'sd-152, 12'sd1815, 13'sd2896}, {12'sd-1083, 9'sd-193, 12'sd-1636}, {12'sd-1129, 13'sd2054, 8'sd79}},
{{12'sd1059, 11'sd832, 12'sd1612}, {13'sd-2413, 12'sd1549, 13'sd2259}, {11'sd-879, 12'sd-1506, 12'sd1572}},
{{12'sd1995, 8'sd107, 13'sd2090}, {13'sd-2387, 9'sd156, 13'sd2655}, {13'sd-2738, 10'sd334, 11'sd628}},
{{12'sd-1181, 13'sd2330, 9'sd-203}, {13'sd2280, 12'sd-1721, 11'sd-941}, {12'sd-1515, 13'sd-2452, 9'sd-192}},
{{12'sd-2012, 12'sd-1410, 10'sd491}, {11'sd-611, 9'sd-207, 11'sd780}, {13'sd2564, 13'sd-2611, 10'sd494}},
{{13'sd2834, 7'sd41, 11'sd730}, {11'sd-797, 12'sd1705, 12'sd-1486}, {13'sd-2096, 13'sd2494, 13'sd2606}},
{{13'sd-2452, 12'sd1419, 12'sd-1419}, {9'sd-212, 13'sd-2812, 13'sd2155}, {8'sd-96, 10'sd339, 13'sd-2920}},
{{9'sd-176, 13'sd2627, 12'sd-1486}, {13'sd2603, 13'sd-2117, 12'sd-1476}, {11'sd528, 10'sd-348, 12'sd1965}},
{{12'sd-1367, 12'sd-1984, 11'sd773}, {9'sd175, 12'sd1953, 12'sd1302}, {7'sd44, 13'sd-2112, 12'sd-2045}},
{{12'sd-1721, 13'sd-2581, 8'sd110}, {12'sd-1503, 9'sd-239, 12'sd1544}, {11'sd1003, 12'sd1563, 10'sd-363}},
{{12'sd2003, 12'sd1425, 13'sd2633}, {8'sd107, 9'sd212, 11'sd760}, {13'sd2097, 11'sd906, 12'sd-1685}},
{{13'sd2632, 8'sd-123, 7'sd57}, {12'sd2046, 13'sd-2343, 10'sd-361}, {13'sd-2625, 13'sd-2230, 13'sd2191}},
{{12'sd-1557, 12'sd2016, 13'sd-3039}, {13'sd2968, 13'sd2084, 10'sd332}, {13'sd2201, 12'sd1610, 13'sd-2748}},
{{13'sd2092, 11'sd-557, 13'sd2692}, {12'sd1636, 13'sd3211, 12'sd1418}, {12'sd-1613, 11'sd651, 11'sd-723}},
{{10'sd478, 12'sd1802, 13'sd2055}, {12'sd-1525, 12'sd1402, 10'sd-340}, {13'sd2286, 13'sd-2298, 13'sd2056}},
{{12'sd-1840, 6'sd-22, 12'sd-1251}, {12'sd1565, 12'sd-1168, 13'sd2289}, {13'sd-2751, 13'sd-2866, 12'sd-1639}},
{{10'sd-406, 11'sd848, 12'sd-1086}, {11'sd-918, 13'sd2136, 8'sd73}, {13'sd3235, 13'sd2467, 11'sd-984}},
{{11'sd-751, 12'sd-1155, 12'sd1083}, {10'sd486, 10'sd-370, 12'sd-1926}, {12'sd1157, 12'sd1681, 13'sd2070}},
{{13'sd-2509, 13'sd-3368, 13'sd-3690}, {12'sd1286, 12'sd-1132, 12'sd-1123}, {13'sd2859, 12'sd-1922, 8'sd97}},
{{12'sd1166, 13'sd-2327, 12'sd-1976}, {13'sd-2240, 13'sd-2352, 11'sd692}, {11'sd831, 11'sd926, 13'sd2585}},
{{12'sd1313, 13'sd-2336, 12'sd-1405}, {8'sd103, 8'sd-95, 10'sd-465}, {12'sd1366, 13'sd2648, 11'sd-895}},
{{10'sd493, 10'sd259, 13'sd-2937}, {13'sd-2329, 11'sd982, 12'sd1629}, {8'sd93, 12'sd-1495, 12'sd-1637}},
{{10'sd-366, 10'sd-420, 11'sd-996}, {12'sd-1913, 12'sd1553, 12'sd1039}, {13'sd-2598, 11'sd-536, 12'sd-1447}},
{{12'sd-1716, 8'sd-99, 12'sd1288}, {12'sd-1037, 12'sd1101, 13'sd2596}, {12'sd1115, 13'sd-2062, 13'sd2202}},
{{9'sd-146, 12'sd-1232, 13'sd2197}, {10'sd-336, 11'sd-636, 9'sd-161}, {12'sd1058, 13'sd-2127, 12'sd1441}},
{{13'sd2589, 7'sd-42, 13'sd-2259}, {13'sd2426, 12'sd-1045, 12'sd1843}, {12'sd-1709, 12'sd1898, 12'sd-1739}},
{{13'sd-2225, 13'sd2167, 11'sd980}, {13'sd-4048, 11'sd955, 11'sd585}, {12'sd-1243, 11'sd-950, 12'sd-1148}},
{{11'sd915, 12'sd-1683, 13'sd2926}, {12'sd1256, 10'sd297, 11'sd-546}, {12'sd-1297, 13'sd2491, 12'sd-1812}},
{{11'sd992, 8'sd-97, 11'sd-962}, {13'sd2702, 12'sd-1593, 13'sd2181}, {10'sd262, 12'sd-1407, 13'sd-2930}},
{{12'sd1588, 10'sd405, 13'sd-2998}, {13'sd2544, 11'sd933, 12'sd1871}, {11'sd-751, 12'sd-1284, 12'sd2036}},
{{9'sd245, 12'sd-1068, 13'sd2490}, {11'sd-894, 10'sd-313, 13'sd2735}, {12'sd-1488, 9'sd182, 10'sd388}},
{{4'sd6, 10'sd477, 9'sd-182}, {12'sd-1387, 12'sd1731, 10'sd-409}, {12'sd-1535, 12'sd1234, 13'sd-2244}},
{{12'sd1349, 12'sd1980, 11'sd603}, {12'sd1973, 13'sd2263, 7'sd-36}, {13'sd2585, 9'sd-139, 13'sd-2672}},
{{12'sd-1200, 13'sd-2800, 11'sd910}, {12'sd1640, 12'sd2032, 12'sd1462}, {11'sd826, 8'sd-87, 12'sd-1041}}},
{
{{12'sd-1188, 12'sd1389, 13'sd-2199}, {12'sd1745, 12'sd1866, 12'sd-1695}, {11'sd-770, 12'sd-1386, 13'sd-2069}},
{{10'sd-437, 10'sd411, 12'sd-1536}, {13'sd2153, 10'sd290, 12'sd-1962}, {12'sd1429, 11'sd-760, 13'sd-2361}},
{{12'sd1730, 8'sd-89, 12'sd1829}, {12'sd-1442, 12'sd1583, 12'sd2032}, {13'sd2065, 13'sd2593, 13'sd-2319}},
{{12'sd1388, 12'sd1809, 12'sd-1150}, {13'sd2950, 11'sd-809, 7'sd-40}, {12'sd-1787, 12'sd-1666, 6'sd-17}},
{{13'sd2317, 8'sd-86, 13'sd2176}, {10'sd325, 13'sd2542, 12'sd-1384}, {12'sd1284, 10'sd449, 12'sd1198}},
{{13'sd-2873, 13'sd-3499, 14'sd-4650}, {13'sd2251, 12'sd1789, 13'sd-2582}, {12'sd1482, 13'sd-2658, 13'sd-3676}},
{{13'sd3670, 12'sd1808, 12'sd-1873}, {12'sd1986, 11'sd907, 12'sd1276}, {12'sd1318, 13'sd2371, 12'sd-1103}},
{{12'sd1761, 13'sd2472, 11'sd795}, {12'sd-1158, 11'sd-627, 13'sd-2475}, {12'sd1764, 8'sd103, 8'sd-109}},
{{11'sd924, 13'sd2459, 13'sd2182}, {11'sd-853, 13'sd2333, 12'sd-1857}, {12'sd1536, 11'sd-816, 12'sd1535}},
{{12'sd2037, 11'sd564, 12'sd-1668}, {8'sd-94, 13'sd-2364, 12'sd1311}, {12'sd-1896, 11'sd-718, 12'sd2010}},
{{12'sd-1084, 11'sd938, 12'sd1202}, {10'sd-369, 11'sd718, 9'sd-159}, {12'sd1232, 10'sd385, 12'sd-1754}},
{{12'sd-1536, 11'sd521, 13'sd-2712}, {11'sd-811, 11'sd-960, 12'sd1088}, {13'sd2312, 12'sd-1268, 11'sd938}},
{{13'sd-2243, 12'sd1575, 12'sd1509}, {12'sd-1317, 13'sd-2627, 11'sd-832}, {12'sd-1646, 12'sd1651, 12'sd-2024}},
{{11'sd-754, 11'sd1007, 11'sd-620}, {10'sd351, 12'sd-1460, 11'sd648}, {13'sd2751, 11'sd-698, 12'sd1802}},
{{11'sd-845, 8'sd-97, 13'sd3791}, {11'sd746, 14'sd4868, 11'sd521}, {13'sd3309, 8'sd93, 14'sd4168}},
{{12'sd-1508, 12'sd-1072, 12'sd1058}, {12'sd-1083, 13'sd-2409, 12'sd-1670}, {12'sd1039, 11'sd925, 12'sd1124}},
{{11'sd819, 12'sd1667, 13'sd-2465}, {13'sd-2911, 13'sd-2463, 9'sd-240}, {10'sd482, 11'sd864, 13'sd2495}},
{{12'sd1241, 12'sd1174, 12'sd-1774}, {12'sd1621, 13'sd2335, 12'sd-1391}, {12'sd-1076, 6'sd-29, 11'sd-817}},
{{8'sd93, 12'sd-1180, 9'sd236}, {12'sd-1431, 12'sd2004, 9'sd-217}, {9'sd-134, 12'sd2043, 13'sd2256}},
{{12'sd-1912, 10'sd420, 12'sd-1499}, {12'sd1349, 12'sd-1864, 10'sd-276}, {13'sd-2350, 13'sd2397, 12'sd1313}},
{{12'sd1381, 13'sd-2562, 12'sd1509}, {12'sd1455, 13'sd-2132, 10'sd419}, {12'sd1403, 11'sd868, 13'sd-2146}},
{{8'sd-80, 7'sd60, 12'sd-1450}, {12'sd-1588, 13'sd2200, 11'sd956}, {12'sd1919, 8'sd108, 12'sd-1660}},
{{13'sd-2388, 12'sd1316, 13'sd2119}, {12'sd1904, 12'sd-1171, 12'sd1875}, {13'sd-2740, 13'sd-2073, 11'sd-645}},
{{10'sd443, 11'sd-864, 12'sd-1585}, {10'sd-287, 11'sd-990, 13'sd-2256}, {12'sd-1040, 13'sd-2255, 13'sd-2084}},
{{13'sd-2149, 11'sd699, 13'sd2329}, {12'sd-1678, 11'sd-858, 13'sd2770}, {13'sd2493, 12'sd-1648, 12'sd1349}},
{{13'sd-2392, 11'sd-746, 12'sd-1262}, {12'sd1220, 11'sd898, 12'sd1702}, {12'sd-1084, 11'sd-668, 11'sd715}},
{{12'sd1877, 10'sd477, 12'sd1504}, {13'sd2132, 12'sd1463, 12'sd-1882}, {13'sd3911, 12'sd1638, 13'sd-2119}},
{{11'sd-655, 11'sd-753, 13'sd-2444}, {9'sd136, 12'sd1102, 11'sd827}, {12'sd1389, 10'sd-281, 11'sd-693}},
{{11'sd-629, 12'sd-1944, 10'sd464}, {12'sd-1397, 12'sd1375, 7'sd51}, {13'sd-2139, 12'sd1681, 11'sd842}},
{{11'sd-725, 6'sd-25, 13'sd2476}, {12'sd1305, 10'sd-304, 12'sd1154}, {13'sd2616, 12'sd1812, 13'sd2602}},
{{12'sd1902, 12'sd1024, 12'sd-1551}, {10'sd487, 10'sd307, 11'sd1001}, {12'sd1099, 11'sd1016, 11'sd888}},
{{12'sd-1654, 12'sd1916, 12'sd-1325}, {13'sd-2346, 12'sd1537, 12'sd-1734}, {13'sd-2994, 13'sd-2251, 13'sd2144}},
{{7'sd-61, 12'sd1124, 13'sd2128}, {12'sd-1377, 12'sd1685, 12'sd-1056}, {12'sd-1689, 13'sd-2125, 12'sd-1329}},
{{12'sd1173, 12'sd-1077, 11'sd696}, {11'sd-972, 13'sd2372, 12'sd1632}, {13'sd2096, 10'sd295, 13'sd2804}},
{{5'sd9, 12'sd-1153, 11'sd-658}, {12'sd1730, 13'sd-2111, 11'sd-588}, {12'sd-1126, 11'sd782, 13'sd2975}},
{{12'sd2019, 12'sd-1695, 11'sd796}, {13'sd-2180, 10'sd294, 13'sd2445}, {13'sd2280, 7'sd37, 11'sd831}},
{{13'sd-3176, 13'sd-3599, 10'sd-413}, {11'sd668, 11'sd-670, 11'sd-892}, {12'sd2014, 13'sd-2257, 13'sd2389}},
{{10'sd-436, 11'sd-742, 12'sd1200}, {12'sd1369, 13'sd-2101, 12'sd1790}, {11'sd798, 11'sd-818, 12'sd1050}},
{{12'sd1303, 12'sd1476, 13'sd-2422}, {12'sd1770, 13'sd2374, 11'sd-736}, {11'sd550, 12'sd1519, 12'sd-1683}},
{{11'sd997, 12'sd-1842, 12'sd-1893}, {12'sd-1882, 13'sd-2642, 12'sd-1359}, {7'sd39, 10'sd448, 12'sd1184}},
{{10'sd306, 10'sd277, 8'sd-124}, {9'sd-141, 11'sd-762, 11'sd-830}, {11'sd992, 13'sd-2142, 12'sd1517}},
{{13'sd-2343, 11'sd-686, 12'sd1266}, {11'sd-572, 12'sd-1904, 13'sd-2765}, {12'sd1538, 11'sd907, 12'sd1639}},
{{12'sd1482, 10'sd499, 12'sd1825}, {3'sd-3, 12'sd-1113, 12'sd1569}, {11'sd-949, 12'sd1379, 8'sd-98}},
{{10'sd390, 13'sd-2334, 13'sd-3206}, {12'sd1433, 12'sd1358, 14'sd-4144}, {10'sd270, 12'sd1426, 12'sd-1193}},
{{13'sd2550, 10'sd482, 12'sd1881}, {11'sd-783, 11'sd-586, 12'sd1151}, {12'sd-1856, 12'sd-1409, 13'sd-2577}},
{{11'sd-972, 11'sd-573, 13'sd2148}, {13'sd2366, 12'sd1596, 10'sd-472}, {11'sd607, 10'sd313, 11'sd-880}},
{{11'sd-886, 11'sd746, 11'sd-753}, {10'sd443, 12'sd-1646, 10'sd-270}, {11'sd-896, 12'sd1845, 13'sd-2648}},
{{13'sd2222, 13'sd2848, 10'sd-294}, {12'sd1506, 13'sd3023, 12'sd1981}, {12'sd1043, 11'sd899, 10'sd-411}},
{{13'sd-2240, 7'sd32, 12'sd1551}, {13'sd3181, 13'sd2888, 13'sd-2529}, {12'sd1910, 11'sd933, 12'sd1793}},
{{12'sd-1828, 11'sd1001, 13'sd-2130}, {13'sd-3868, 13'sd-3700, 13'sd2619}, {11'sd-1018, 10'sd405, 11'sd603}},
{{12'sd1056, 7'sd42, 12'sd-1276}, {13'sd-2630, 12'sd-1752, 11'sd-1016}, {9'sd-215, 11'sd-519, 13'sd3061}},
{{13'sd-2106, 12'sd1573, 12'sd-1188}, {13'sd-2872, 10'sd361, 13'sd-2856}, {11'sd817, 12'sd-1335, 9'sd224}},
{{10'sd296, 12'sd1766, 12'sd1029}, {10'sd411, 13'sd2812, 11'sd954}, {9'sd-229, 11'sd-733, 12'sd1641}},
{{13'sd2461, 13'sd2694, 13'sd-2194}, {10'sd-372, 11'sd-564, 9'sd135}, {13'sd-2165, 13'sd-2473, 10'sd475}},
{{13'sd3892, 11'sd-583, 9'sd-230}, {13'sd2728, 11'sd917, 11'sd942}, {12'sd-1418, 13'sd-2161, 11'sd-621}},
{{11'sd-908, 13'sd-3020, 13'sd2277}, {12'sd-1695, 8'sd65, 13'sd2380}, {12'sd-1179, 13'sd-2085, 13'sd2252}},
{{12'sd1660, 12'sd1229, 13'sd3011}, {12'sd-2031, 12'sd-1766, 13'sd2664}, {13'sd2690, 13'sd2845, 12'sd-1697}},
{{12'sd1354, 13'sd2074, 11'sd-799}, {13'sd2313, 13'sd-2297, 13'sd2327}, {13'sd-2514, 11'sd1012, 12'sd1042}},
{{13'sd2403, 11'sd-1006, 12'sd-1667}, {11'sd-829, 10'sd499, 12'sd-1806}, {7'sd50, 12'sd1460, 13'sd-2671}},
{{12'sd-1813, 12'sd1284, 10'sd-308}, {11'sd932, 12'sd1430, 12'sd1077}, {13'sd3032, 12'sd1102, 11'sd-723}},
{{10'sd257, 13'sd-2471, 9'sd210}, {13'sd-2428, 12'sd1983, 11'sd-708}, {12'sd-1834, 7'sd43, 12'sd1427}},
{{8'sd-95, 12'sd1524, 12'sd-1292}, {13'sd-2665, 11'sd-770, 13'sd-2382}, {8'sd-96, 11'sd-521, 12'sd1216}},
{{11'sd-629, 4'sd-6, 10'sd-388}, {13'sd-2378, 11'sd695, 12'sd-1111}, {12'sd1521, 13'sd-2061, 10'sd-454}},
{{13'sd-2658, 13'sd-2101, 12'sd1695}, {11'sd545, 10'sd-264, 12'sd1184}, {12'sd1753, 11'sd-714, 12'sd-1222}}},
{
{{9'sd-223, 12'sd-1370, 13'sd-2186}, {13'sd2281, 13'sd2489, 11'sd-970}, {13'sd2720, 11'sd530, 12'sd-1430}},
{{10'sd300, 11'sd-748, 12'sd1609}, {11'sd807, 12'sd1340, 7'sd34}, {9'sd161, 9'sd219, 10'sd305}},
{{13'sd4037, 13'sd2676, 10'sd354}, {12'sd-1190, 11'sd870, 9'sd-199}, {10'sd416, 12'sd1726, 11'sd-951}},
{{11'sd602, 10'sd-341, 10'sd440}, {12'sd-1760, 12'sd-1743, 12'sd1236}, {12'sd-1859, 12'sd-1169, 12'sd-1341}},
{{11'sd672, 11'sd-1005, 13'sd2265}, {12'sd1091, 12'sd1756, 12'sd-1380}, {10'sd256, 7'sd-53, 12'sd-1701}},
{{13'sd-3648, 10'sd404, 13'sd2272}, {12'sd-1932, 10'sd325, 12'sd1554}, {13'sd-3540, 10'sd317, 14'sd-4542}},
{{13'sd-2513, 12'sd-1316, 12'sd-1105}, {14'sd-5169, 11'sd673, 10'sd-425}, {12'sd-1730, 13'sd-2129, 13'sd-2132}},
{{13'sd-2935, 9'sd154, 11'sd768}, {13'sd-2243, 12'sd-1371, 12'sd-1364}, {11'sd-602, 12'sd1263, 12'sd-1583}},
{{11'sd-829, 9'sd239, 13'sd-2588}, {13'sd-2201, 8'sd-79, 13'sd2198}, {9'sd245, 10'sd473, 12'sd-1650}},
{{12'sd-1082, 11'sd-677, 12'sd-1283}, {12'sd-1921, 11'sd-937, 12'sd-1823}, {10'sd-330, 12'sd-1635, 13'sd-2320}},
{{14'sd4651, 13'sd3701, 13'sd2921}, {13'sd2223, 10'sd497, 10'sd361}, {10'sd412, 11'sd-529, 13'sd3114}},
{{11'sd548, 13'sd2941, 12'sd-1861}, {12'sd-1151, 11'sd-656, 8'sd86}, {13'sd3046, 13'sd-2050, 11'sd-828}},
{{11'sd813, 13'sd-3096, 12'sd1584}, {12'sd-1200, 13'sd-2839, 12'sd-1253}, {7'sd-63, 13'sd-2468, 12'sd-1927}},
{{11'sd-770, 12'sd1440, 13'sd2340}, {12'sd1471, 10'sd410, 13'sd2519}, {13'sd2554, 12'sd1146, 12'sd1065}},
{{10'sd462, 12'sd-1385, 12'sd-1240}, {13'sd-2993, 14'sd-5479, 12'sd-1920}, {14'sd-4350, 14'sd-4487, 14'sd-4127}},
{{13'sd3259, 12'sd-1266, 13'sd-2672}, {11'sd-998, 12'sd-1076, 12'sd1277}, {9'sd171, 13'sd-2340, 11'sd1017}},
{{12'sd-1444, 12'sd-1208, 13'sd-2624}, {12'sd1689, 13'sd2723, 11'sd-864}, {12'sd1891, 11'sd707, 13'sd2579}},
{{12'sd-1881, 11'sd998, 12'sd1606}, {13'sd2134, 11'sd-528, 13'sd-2479}, {11'sd598, 8'sd-126, 14'sd-4515}},
{{9'sd226, 12'sd1106, 13'sd-3196}, {13'sd2348, 13'sd-2645, 12'sd-2002}, {5'sd-12, 13'sd-2940, 12'sd-1950}},
{{13'sd-2972, 13'sd-2652, 12'sd-1031}, {12'sd-1230, 13'sd2290, 11'sd-828}, {12'sd-1091, 13'sd-2580, 11'sd767}},
{{13'sd-3188, 11'sd-816, 12'sd-1420}, {12'sd-1491, 12'sd2007, 12'sd-1221}, {12'sd-1952, 9'sd-218, 13'sd-2136}},
{{12'sd1984, 6'sd16, 13'sd2332}, {10'sd-330, 12'sd-1189, 13'sd2256}, {12'sd1335, 12'sd-1173, 12'sd-1631}},
{{11'sd-731, 9'sd241, 11'sd-776}, {12'sd-1316, 13'sd2464, 13'sd2295}, {13'sd3312, 6'sd-30, 11'sd729}},
{{10'sd335, 13'sd-2989, 12'sd-1498}, {11'sd953, 11'sd-610, 12'sd-1539}, {12'sd1477, 12'sd-1236, 12'sd1166}},
{{10'sd257, 13'sd2429, 12'sd1550}, {12'sd1208, 12'sd-1657, 13'sd2541}, {12'sd1594, 11'sd-834, 11'sd918}},
{{11'sd-772, 9'sd-214, 12'sd-2007}, {10'sd-399, 12'sd-1065, 10'sd356}, {13'sd2178, 11'sd-706, 13'sd-2796}},
{{13'sd3455, 14'sd4831, 13'sd2340}, {14'sd5403, 12'sd1692, 10'sd451}, {13'sd-2379, 12'sd-1162, 8'sd104}},
{{13'sd-2456, 12'sd-2014, 13'sd2465}, {9'sd215, 12'sd-1395, 13'sd-2101}, {11'sd693, 13'sd-2516, 14'sd-4141}},
{{13'sd3009, 12'sd-1787, 12'sd1712}, {11'sd1017, 11'sd728, 11'sd-850}, {12'sd1407, 11'sd-702, 13'sd3290}},
{{13'sd-2486, 9'sd-135, 13'sd2060}, {11'sd948, 10'sd-418, 13'sd2739}, {10'sd-367, 12'sd1855, 12'sd1253}},
{{12'sd-1476, 9'sd215, 11'sd675}, {13'sd-2383, 13'sd2818, 12'sd1514}, {12'sd1290, 13'sd2468, 13'sd2284}},
{{10'sd296, 12'sd1642, 8'sd92}, {13'sd2556, 10'sd-472, 11'sd-726}, {13'sd2170, 12'sd1675, 13'sd2160}},
{{9'sd-182, 12'sd-1751, 13'sd-2064}, {12'sd1900, 8'sd71, 1'sd0}, {13'sd-2118, 12'sd-1328, 13'sd2437}},
{{13'sd2607, 9'sd155, 7'sd48}, {12'sd1114, 13'sd-2889, 13'sd2418}, {11'sd-740, 13'sd-3343, 13'sd-2766}},
{{13'sd-2991, 11'sd733, 12'sd-1191}, {9'sd-128, 11'sd562, 12'sd1536}, {8'sd-66, 11'sd685, 13'sd2494}},
{{12'sd-1200, 11'sd-1004, 9'sd-241}, {12'sd1135, 7'sd48, 10'sd-435}, {11'sd651, 12'sd-1433, 10'sd300}},
{{13'sd-3452, 12'sd1582, 10'sd-378}, {13'sd-2989, 12'sd-1839, 11'sd-639}, {14'sd-6263, 11'sd866, 13'sd2734}},
{{12'sd-1613, 12'sd-1974, 12'sd1113}, {11'sd-816, 11'sd-689, 13'sd-2328}, {13'sd-3488, 11'sd-746, 14'sd-4193}},
{{12'sd-1996, 10'sd274, 11'sd799}, {9'sd-189, 11'sd649, 12'sd1631}, {10'sd298, 13'sd2401, 11'sd562}},
{{12'sd-1150, 13'sd-2523, 11'sd-680}, {13'sd2372, 13'sd-2461, 12'sd-1050}, {12'sd1706, 12'sd-1686, 12'sd-1287}},
{{13'sd-3105, 9'sd-210, 11'sd800}, {13'sd-2472, 10'sd-342, 13'sd-2100}, {14'sd-7275, 14'sd-4272, 14'sd-4316}},
{{13'sd3214, 12'sd1448, 12'sd1207}, {13'sd3121, 10'sd-479, 11'sd-947}, {10'sd505, 13'sd3112, 13'sd2778}},
{{13'sd3633, 13'sd2980, 13'sd2233}, {10'sd305, 11'sd-768, 12'sd1228}, {13'sd3325, 9'sd224, 11'sd-751}},
{{15'sd12812, 14'sd6715, 15'sd12194}, {15'sd9609, 14'sd4596, 14'sd7195}, {14'sd7994, 14'sd5117, 13'sd3307}},
{{10'sd-369, 7'sd35, 11'sd647}, {4'sd6, 13'sd-2450, 11'sd790}, {12'sd-1826, 13'sd-2654, 13'sd-2882}},
{{13'sd-2570, 12'sd1835, 13'sd2168}, {11'sd-571, 12'sd2014, 12'sd-1453}, {12'sd1754, 13'sd2244, 10'sd-441}},
{{9'sd243, 11'sd-563, 11'sd936}, {11'sd656, 11'sd708, 11'sd718}, {13'sd-3629, 13'sd-2181, 12'sd1070}},
{{11'sd965, 12'sd-1394, 9'sd165}, {11'sd-746, 11'sd-543, 6'sd-22}, {12'sd-1149, 13'sd-2372, 13'sd2572}},
{{12'sd1414, 13'sd4006, 13'sd3608}, {6'sd23, 13'sd2273, 11'sd-575}, {13'sd-2836, 10'sd336, 13'sd2787}},
{{9'sd232, 13'sd-3009, 13'sd-3271}, {12'sd1408, 12'sd1186, 13'sd-2612}, {12'sd1324, 11'sd-868, 12'sd1267}},
{{13'sd-3462, 10'sd-297, 12'sd-1996}, {12'sd-2002, 13'sd2910, 11'sd-754}, {11'sd876, 12'sd-1115, 13'sd-2744}},
{{11'sd-858, 11'sd872, 9'sd-176}, {13'sd2677, 11'sd-592, 13'sd-2163}, {14'sd4768, 11'sd-675, 12'sd-1519}},
{{12'sd-1937, 11'sd562, 12'sd-1532}, {12'sd-1446, 12'sd1233, 12'sd-1723}, {13'sd2526, 12'sd-1406, 11'sd689}},
{{13'sd2484, 13'sd-2340, 13'sd2380}, {11'sd-599, 9'sd254, 11'sd-598}, {12'sd1859, 12'sd1281, 12'sd1028}},
{{13'sd-3940, 12'sd-1730, 8'sd-84}, {12'sd1168, 13'sd-3653, 12'sd-1663}, {13'sd-3024, 8'sd-81, 13'sd-3599}},
{{13'sd-3392, 12'sd1099, 11'sd803}, {12'sd-1261, 7'sd37, 12'sd1517}, {12'sd-1279, 13'sd2664, 12'sd-1633}},
{{12'sd-1574, 11'sd629, 10'sd495}, {13'sd-2297, 13'sd-3254, 13'sd-3998}, {14'sd7159, 13'sd3875, 13'sd2154}},
{{12'sd-1120, 12'sd1939, 10'sd-463}, {13'sd-2126, 12'sd-1944, 10'sd506}, {12'sd-1420, 13'sd-2450, 11'sd873}},
{{13'sd2609, 10'sd424, 13'sd2726}, {11'sd917, 13'sd-2864, 12'sd1308}, {9'sd-129, 13'sd-2201, 12'sd-1259}},
{{10'sd-392, 13'sd-2291, 12'sd1351}, {12'sd-1418, 13'sd2337, 12'sd1382}, {13'sd-3775, 14'sd-4934, 12'sd-1293}},
{{12'sd-1749, 8'sd-126, 11'sd-941}, {12'sd1430, 13'sd-2760, 13'sd2213}, {13'sd-2920, 9'sd-189, 12'sd1988}},
{{9'sd231, 10'sd299, 12'sd-1859}, {13'sd-2476, 12'sd-1301, 8'sd-116}, {11'sd653, 10'sd-427, 13'sd2353}},
{{13'sd2070, 10'sd-456, 12'sd-1260}, {12'sd-1977, 12'sd1661, 11'sd650}, {11'sd965, 12'sd-1341, 13'sd2916}},
{{12'sd1678, 13'sd3001, 11'sd924}, {13'sd3777, 11'sd624, 12'sd1946}, {12'sd-1523, 12'sd-1779, 13'sd3334}}},
{
{{13'sd-2173, 13'sd-2308, 12'sd1638}, {12'sd-1717, 13'sd2730, 12'sd1333}, {9'sd238, 12'sd1030, 13'sd-2307}},
{{11'sd883, 12'sd1613, 13'sd2113}, {12'sd-1427, 11'sd-795, 12'sd-1787}, {11'sd-632, 12'sd2005, 12'sd-2018}},
{{13'sd2585, 12'sd-1996, 12'sd-1664}, {13'sd-2362, 13'sd2183, 12'sd1071}, {12'sd-1966, 13'sd-2845, 11'sd-929}},
{{12'sd2031, 12'sd1046, 13'sd2486}, {12'sd-1836, 13'sd-2747, 9'sd161}, {12'sd-1203, 12'sd-1435, 13'sd-2148}},
{{12'sd-1830, 11'sd871, 12'sd1221}, {12'sd-2037, 11'sd-653, 13'sd-3179}, {12'sd-1062, 8'sd106, 13'sd-3713}},
{{12'sd1540, 11'sd-800, 12'sd1461}, {7'sd60, 13'sd-2325, 13'sd2136}, {11'sd-548, 12'sd1773, 12'sd1643}},
{{11'sd753, 13'sd-2452, 13'sd-2433}, {13'sd-2892, 6'sd-17, 13'sd-2191}, {11'sd-930, 13'sd-2768, 8'sd77}},
{{12'sd-1720, 12'sd1451, 11'sd-622}, {12'sd1337, 12'sd1675, 11'sd-932}, {12'sd-1619, 10'sd-474, 10'sd-396}},
{{11'sd885, 8'sd-83, 11'sd-649}, {8'sd102, 12'sd2012, 12'sd1024}, {12'sd1887, 12'sd1642, 13'sd2579}},
{{12'sd-1804, 12'sd1407, 11'sd893}, {12'sd-1958, 12'sd-1904, 13'sd-2834}, {11'sd-826, 10'sd362, 9'sd-212}},
{{12'sd-1205, 13'sd-2739, 9'sd-222}, {12'sd-1532, 11'sd-680, 11'sd-577}, {12'sd-1670, 12'sd-1091, 12'sd-1639}},
{{12'sd-1955, 12'sd-2029, 12'sd1563}, {12'sd-2027, 13'sd2260, 12'sd-1558}, {10'sd-477, 10'sd-282, 11'sd-889}},
{{12'sd-1789, 11'sd1005, 10'sd-296}, {12'sd-2001, 12'sd-1831, 12'sd1971}, {13'sd2133, 13'sd2347, 11'sd-578}},
{{13'sd-2380, 12'sd-1416, 13'sd-2733}, {12'sd-1581, 10'sd498, 12'sd1108}, {13'sd-2152, 12'sd1361, 13'sd-2467}},
{{11'sd739, 10'sd264, 13'sd-3353}, {12'sd-1914, 5'sd-14, 13'sd-2948}, {12'sd-1315, 9'sd179, 13'sd-2365}},
{{13'sd-2695, 10'sd-330, 11'sd890}, {12'sd1510, 11'sd571, 11'sd-615}, {11'sd-734, 12'sd-1744, 12'sd1323}},
{{11'sd-919, 11'sd690, 9'sd-148}, {12'sd1444, 13'sd2371, 11'sd-855}, {10'sd478, 12'sd-1053, 12'sd-1238}},
{{10'sd364, 12'sd-1918, 12'sd-1862}, {12'sd-1078, 12'sd-1807, 12'sd1597}, {10'sd406, 12'sd-1956, 9'sd-232}},
{{12'sd-1404, 13'sd2360, 11'sd957}, {11'sd942, 13'sd-2417, 13'sd-2615}, {13'sd2631, 11'sd-912, 13'sd-2406}},
{{12'sd-1335, 13'sd2259, 11'sd-543}, {13'sd2268, 11'sd-582, 10'sd362}, {12'sd1296, 11'sd586, 12'sd-1660}},
{{12'sd1202, 13'sd2702, 11'sd614}, {12'sd-1674, 12'sd1577, 12'sd-1488}, {12'sd1389, 7'sd49, 10'sd-302}},
{{13'sd2475, 13'sd2499, 12'sd1153}, {7'sd-63, 12'sd1185, 12'sd1728}, {13'sd2337, 13'sd2494, 12'sd1271}},
{{10'sd295, 12'sd-1320, 13'sd2466}, {9'sd208, 13'sd2149, 13'sd2457}, {12'sd1089, 11'sd-560, 12'sd1431}},
{{13'sd-2601, 13'sd-2523, 13'sd2179}, {13'sd2178, 10'sd-437, 11'sd-982}, {13'sd2560, 12'sd1508, 12'sd-1310}},
{{12'sd1977, 13'sd-2712, 13'sd-2814}, {9'sd170, 12'sd1111, 13'sd-2720}, {13'sd2535, 11'sd-699, 12'sd1108}},
{{13'sd-2401, 8'sd71, 12'sd-1459}, {11'sd-586, 13'sd2131, 11'sd1004}, {13'sd-2564, 11'sd780, 12'sd-1720}},
{{13'sd-2147, 13'sd-3287, 13'sd-3090}, {14'sd-4750, 13'sd-3175, 13'sd-3594}, {8'sd-73, 13'sd-3224, 12'sd1135}},
{{12'sd-1553, 13'sd-2295, 10'sd330}, {12'sd-1612, 11'sd948, 11'sd-854}, {11'sd773, 10'sd-449, 12'sd1737}},
{{12'sd-1631, 12'sd1822, 11'sd991}, {11'sd1021, 10'sd-424, 12'sd-1239}, {13'sd-2611, 11'sd707, 11'sd-838}},
{{13'sd-2843, 12'sd-1666, 13'sd-2524}, {13'sd-3358, 11'sd782, 12'sd-1175}, {12'sd1298, 12'sd1470, 12'sd-1666}},
{{12'sd-1898, 12'sd1139, 12'sd1333}, {12'sd-1227, 10'sd-405, 13'sd2247}, {11'sd891, 11'sd962, 13'sd2174}},
{{11'sd549, 13'sd2628, 13'sd-2670}, {11'sd-990, 5'sd-8, 12'sd-1564}, {12'sd1064, 9'sd160, 13'sd-2209}},
{{9'sd-213, 13'sd2197, 12'sd-1610}, {10'sd-389, 11'sd-985, 11'sd-783}, {11'sd582, 12'sd1219, 12'sd2029}},
{{11'sd782, 12'sd1502, 11'sd679}, {11'sd-729, 12'sd1038, 9'sd169}, {12'sd1135, 10'sd305, 12'sd1586}},
{{13'sd-2079, 13'sd2465, 10'sd-257}, {13'sd2495, 9'sd-235, 13'sd3058}, {12'sd-1034, 9'sd239, 13'sd2363}},
{{13'sd2410, 13'sd2422, 11'sd-754}, {12'sd1900, 11'sd678, 13'sd-2648}, {11'sd-547, 13'sd2426, 12'sd-1413}},
{{12'sd1060, 6'sd17, 11'sd-737}, {12'sd-1799, 10'sd310, 13'sd3876}, {11'sd698, 9'sd-195, 13'sd2412}},
{{10'sd416, 11'sd-679, 8'sd-70}, {13'sd-2551, 13'sd-2735, 12'sd-1935}, {13'sd-2939, 9'sd-159, 7'sd-34}},
{{13'sd2681, 12'sd1741, 10'sd367}, {13'sd-2837, 12'sd1148, 13'sd-2101}, {13'sd-2831, 11'sd661, 13'sd2627}},
{{9'sd-202, 12'sd-1591, 13'sd-2094}, {11'sd870, 13'sd2275, 12'sd1960}, {12'sd-1855, 10'sd342, 12'sd-1272}},
{{12'sd-1975, 13'sd-2493, 13'sd-2705}, {12'sd1539, 13'sd-3011, 7'sd-35}, {12'sd-1195, 11'sd932, 12'sd-1440}},
{{12'sd1139, 11'sd-889, 13'sd-2176}, {13'sd-2347, 13'sd-2814, 12'sd-1094}, {11'sd762, 12'sd1952, 11'sd722}},
{{13'sd-2653, 10'sd-469, 9'sd-164}, {10'sd330, 12'sd-1595, 13'sd-3020}, {13'sd-2571, 12'sd-1420, 12'sd1154}},
{{10'sd413, 12'sd1812, 12'sd1733}, {13'sd-3916, 11'sd773, 13'sd2926}, {13'sd-3970, 13'sd-3797, 13'sd-3309}},
{{11'sd612, 13'sd-2132, 12'sd-1680}, {12'sd1393, 12'sd1136, 12'sd-1415}, {13'sd-2300, 9'sd138, 13'sd2107}},
{{12'sd-1402, 6'sd17, 8'sd-82}, {12'sd-1825, 12'sd1786, 13'sd2212}, {12'sd1027, 11'sd832, 12'sd1829}},
{{12'sd1353, 13'sd-2170, 12'sd1041}, {12'sd-1076, 13'sd2356, 12'sd-1872}, {11'sd963, 11'sd-832, 11'sd-798}},
{{11'sd760, 11'sd-811, 11'sd721}, {13'sd-2396, 12'sd-1957, 8'sd-89}, {12'sd-1561, 12'sd-1304, 12'sd1185}},
{{12'sd-1549, 12'sd1114, 12'sd-1694}, {12'sd1514, 10'sd-422, 12'sd-1585}, {13'sd-2089, 9'sd-166, 12'sd-1179}},
{{13'sd2063, 11'sd-521, 12'sd-1648}, {13'sd2377, 12'sd1161, 12'sd1138}, {13'sd3741, 12'sd1881, 12'sd1380}},
{{12'sd-2018, 11'sd910, 6'sd30}, {13'sd2464, 11'sd-532, 12'sd-1055}, {12'sd1096, 13'sd-2402, 10'sd340}},
{{11'sd-540, 11'sd684, 12'sd1126}, {12'sd1964, 12'sd1258, 12'sd-1246}, {12'sd-1666, 12'sd-1583, 10'sd-452}},
{{12'sd-1166, 13'sd2890, 12'sd1637}, {12'sd2038, 11'sd-884, 11'sd805}, {12'sd-1669, 11'sd-726, 10'sd337}},
{{13'sd2294, 9'sd-243, 12'sd-1399}, {12'sd1600, 12'sd-1375, 12'sd-1476}, {12'sd-1634, 12'sd-1419, 12'sd-1039}},
{{13'sd-3164, 11'sd-1005, 10'sd478}, {12'sd-1815, 13'sd-3185, 10'sd383}, {13'sd-3059, 13'sd-2206, 9'sd-179}},
{{12'sd-1146, 12'sd1595, 12'sd-1035}, {12'sd-1099, 13'sd2509, 10'sd-288}, {12'sd1580, 12'sd-1732, 9'sd151}},
{{9'sd141, 13'sd-3528, 13'sd-3852}, {12'sd-1881, 12'sd-1927, 13'sd-2562}, {12'sd-1447, 13'sd-3236, 13'sd-2452}},
{{11'sd647, 12'sd1307, 10'sd-408}, {12'sd1985, 10'sd-400, 11'sd-668}, {13'sd-2401, 11'sd-1016, 13'sd2130}},
{{11'sd663, 13'sd-2178, 11'sd-586}, {13'sd-2873, 13'sd-2210, 12'sd-1589}, {12'sd-1960, 13'sd-2923, 12'sd2028}},
{{10'sd-361, 13'sd-2076, 8'sd-124}, {12'sd1298, 13'sd2136, 11'sd853}, {11'sd-653, 10'sd349, 12'sd1208}},
{{12'sd1365, 12'sd1684, 13'sd2733}, {13'sd2174, 12'sd-1953, 10'sd500}, {12'sd1315, 10'sd382, 12'sd-1349}},
{{12'sd-1437, 10'sd-347, 12'sd-2025}, {10'sd-480, 11'sd-549, 12'sd1119}, {13'sd2358, 13'sd2243, 12'sd1470}},
{{12'sd-1232, 11'sd727, 12'sd1303}, {13'sd-2128, 12'sd1037, 11'sd-748}, {11'sd735, 10'sd331, 12'sd-1053}},
{{9'sd138, 12'sd1550, 12'sd-1598}, {10'sd298, 5'sd-14, 12'sd-1163}, {11'sd-928, 10'sd-450, 8'sd118}}},
{
{{11'sd989, 11'sd642, 8'sd113}, {9'sd201, 12'sd2000, 12'sd-1903}, {13'sd2381, 12'sd1994, 10'sd-419}},
{{12'sd1567, 11'sd1007, 12'sd1948}, {13'sd-2130, 9'sd231, 6'sd-19}, {13'sd2829, 13'sd2335, 12'sd-1478}},
{{11'sd690, 5'sd8, 13'sd-2171}, {11'sd616, 13'sd-2869, 10'sd-405}, {13'sd-2381, 12'sd-1810, 11'sd-853}},
{{13'sd-2166, 13'sd2060, 13'sd2500}, {13'sd-2407, 12'sd1247, 11'sd-596}, {13'sd-2824, 13'sd2347, 11'sd-744}},
{{13'sd2152, 11'sd731, 9'sd-237}, {11'sd917, 6'sd-31, 11'sd-866}, {14'sd-4555, 10'sd-261, 13'sd-2147}},
{{11'sd-881, 12'sd-1039, 11'sd-652}, {12'sd-1083, 13'sd2749, 10'sd257}, {10'sd-318, 11'sd-848, 13'sd2451}},
{{12'sd-1211, 11'sd852, 13'sd-2250}, {12'sd1259, 11'sd-786, 13'sd-2371}, {11'sd743, 12'sd-1395, 13'sd-2264}},
{{12'sd-1507, 13'sd2141, 13'sd2123}, {9'sd-157, 13'sd2394, 12'sd-1689}, {11'sd-905, 11'sd-695, 11'sd-538}},
{{10'sd273, 11'sd685, 12'sd-1059}, {11'sd972, 6'sd25, 10'sd391}, {6'sd24, 10'sd431, 12'sd1325}},
{{13'sd-2413, 12'sd-1636, 13'sd-2279}, {12'sd1706, 13'sd-2499, 12'sd-1870}, {12'sd1211, 8'sd80, 11'sd589}},
{{13'sd-2303, 9'sd205, 11'sd-622}, {13'sd-2480, 10'sd-411, 12'sd2038}, {12'sd1081, 12'sd1196, 12'sd-1770}},
{{13'sd2550, 7'sd-53, 12'sd1381}, {9'sd225, 13'sd-2448, 9'sd152}, {12'sd1504, 12'sd-1810, 9'sd-216}},
{{11'sd-872, 11'sd-882, 11'sd-682}, {12'sd1463, 12'sd-1464, 10'sd-257}, {12'sd1834, 10'sd364, 11'sd888}},
{{11'sd791, 13'sd-2427, 12'sd1370}, {10'sd476, 13'sd-2095, 13'sd2153}, {12'sd1507, 13'sd-2445, 12'sd-1379}},
{{8'sd-90, 13'sd-3472, 13'sd-3870}, {11'sd715, 9'sd-198, 12'sd-1768}, {11'sd-580, 12'sd-1923, 14'sd-4278}},
{{13'sd2443, 11'sd755, 13'sd-2515}, {13'sd-2048, 11'sd-944, 13'sd-2620}, {9'sd-195, 8'sd-94, 12'sd1774}},
{{11'sd645, 10'sd-385, 11'sd881}, {13'sd-2293, 12'sd1323, 12'sd-1816}, {12'sd-1656, 13'sd2336, 12'sd1081}},
{{12'sd-1175, 10'sd-475, 12'sd1809}, {11'sd-913, 12'sd-1869, 10'sd472}, {12'sd1577, 12'sd1962, 12'sd-1058}},
{{13'sd2526, 10'sd-471, 13'sd2449}, {9'sd-154, 10'sd-392, 12'sd-1855}, {13'sd2293, 12'sd-1547, 12'sd1239}},
{{12'sd-1686, 11'sd-526, 12'sd1231}, {13'sd2624, 13'sd2888, 9'sd228}, {13'sd2390, 10'sd-405, 12'sd1483}},
{{12'sd1724, 12'sd1361, 13'sd-2134}, {13'sd-2604, 12'sd-1189, 9'sd128}, {13'sd-2711, 13'sd2415, 9'sd138}},
{{11'sd-697, 12'sd-1300, 13'sd2259}, {12'sd-1823, 13'sd2076, 9'sd250}, {10'sd358, 13'sd2481, 13'sd-2230}},
{{12'sd-1560, 13'sd2390, 13'sd2566}, {13'sd-2144, 11'sd591, 10'sd305}, {12'sd-1564, 12'sd1332, 11'sd968}},
{{11'sd-942, 13'sd2563, 10'sd-319}, {11'sd806, 13'sd-2323, 13'sd-2092}, {8'sd-119, 12'sd1561, 13'sd2189}},
{{12'sd1106, 12'sd1823, 13'sd2377}, {12'sd-1073, 11'sd-1019, 12'sd1440}, {13'sd2113, 13'sd2578, 11'sd1004}},
{{12'sd-1947, 13'sd-2338, 12'sd1398}, {13'sd-2815, 9'sd-235, 9'sd-240}, {12'sd-1819, 8'sd102, 9'sd-149}},
{{10'sd-464, 14'sd-4516, 13'sd2161}, {13'sd-2519, 12'sd-1402, 11'sd-929}, {11'sd811, 13'sd-2899, 12'sd1718}},
{{12'sd-1687, 9'sd-179, 7'sd34}, {11'sd-801, 13'sd-3011, 11'sd-531}, {13'sd-2885, 13'sd-2962, 13'sd-2600}},
{{11'sd-553, 12'sd1500, 13'sd-2603}, {12'sd1606, 12'sd1197, 9'sd208}, {12'sd-1928, 13'sd-2273, 9'sd241}},
{{12'sd-1353, 11'sd-754, 13'sd-2609}, {12'sd1920, 13'sd-2431, 11'sd-859}, {11'sd-694, 10'sd389, 10'sd310}},
{{11'sd-557, 10'sd-400, 12'sd-1859}, {11'sd789, 10'sd391, 13'sd-2376}, {13'sd2230, 9'sd-215, 7'sd50}},
{{12'sd1612, 12'sd1353, 11'sd-992}, {13'sd3118, 11'sd743, 12'sd-2007}, {11'sd717, 11'sd722, 11'sd-975}},
{{12'sd1214, 11'sd-669, 12'sd1046}, {9'sd252, 11'sd-682, 13'sd2161}, {10'sd-482, 13'sd2112, 13'sd2374}},
{{12'sd-1378, 12'sd1936, 11'sd-831}, {13'sd2440, 12'sd1901, 11'sd607}, {13'sd2298, 13'sd-2456, 12'sd1912}},
{{12'sd1278, 12'sd1991, 11'sd548}, {9'sd-149, 12'sd1730, 11'sd-726}, {10'sd421, 11'sd962, 12'sd-1291}},
{{12'sd1858, 11'sd607, 13'sd-2159}, {12'sd1827, 12'sd-1689, 11'sd-595}, {8'sd-69, 11'sd813, 13'sd-2415}},
{{13'sd-2077, 11'sd878, 13'sd2588}, {13'sd-2159, 13'sd2672, 11'sd775}, {13'sd2668, 11'sd-896, 13'sd3226}},
{{13'sd-3003, 11'sd-742, 13'sd-2191}, {8'sd73, 11'sd758, 12'sd-1772}, {13'sd-2934, 11'sd-1017, 9'sd183}},
{{11'sd-640, 13'sd-2439, 12'sd-1519}, {13'sd-2071, 9'sd229, 13'sd2480}, {12'sd1439, 11'sd-564, 13'sd-2092}},
{{10'sd-369, 12'sd1503, 13'sd2145}, {12'sd1838, 13'sd-2252, 13'sd2585}, {13'sd2356, 13'sd-2069, 11'sd782}},
{{13'sd-2900, 12'sd1125, 13'sd2116}, {11'sd-766, 10'sd-418, 12'sd1680}, {13'sd2309, 11'sd830, 13'sd-2066}},
{{13'sd2270, 12'sd1615, 12'sd1900}, {9'sd-135, 11'sd652, 12'sd-1468}, {12'sd1343, 12'sd-1821, 12'sd1955}},
{{13'sd-4073, 12'sd-1557, 11'sd618}, {12'sd-1925, 13'sd-3543, 7'sd53}, {13'sd-2303, 12'sd-1611, 13'sd-2593}},
{{12'sd1147, 13'sd-2872, 12'sd-1423}, {10'sd320, 14'sd-4242, 6'sd-20}, {13'sd-2462, 13'sd-4067, 12'sd1195}},
{{13'sd-2797, 12'sd1571, 12'sd-1090}, {13'sd-2854, 12'sd-1961, 7'sd-49}, {12'sd-1789, 12'sd-1444, 12'sd-1216}},
{{12'sd-1928, 13'sd2303, 12'sd1165}, {12'sd-1868, 11'sd-639, 13'sd2290}, {11'sd619, 11'sd-906, 13'sd2643}},
{{11'sd-835, 10'sd-492, 12'sd2039}, {13'sd2904, 12'sd-1894, 11'sd-872}, {8'sd-88, 13'sd2381, 11'sd-685}},
{{13'sd-3717, 13'sd-2143, 12'sd1296}, {13'sd-2853, 12'sd-1604, 13'sd-2386}, {10'sd-301, 11'sd753, 10'sd-412}},
{{12'sd-2033, 13'sd2386, 12'sd-1192}, {11'sd967, 12'sd1212, 12'sd-1423}, {12'sd1701, 13'sd-2360, 11'sd813}},
{{13'sd3689, 12'sd1191, 11'sd-635}, {11'sd-631, 13'sd3020, 10'sd274}, {11'sd-545, 12'sd1915, 11'sd-934}},
{{12'sd-1061, 12'sd-1034, 12'sd-2002}, {11'sd-823, 12'sd-1538, 13'sd-2181}, {12'sd-1119, 12'sd1338, 12'sd-1794}},
{{13'sd2270, 13'sd-2171, 6'sd-19}, {11'sd790, 12'sd-1180, 12'sd1329}, {10'sd-336, 12'sd-1744, 11'sd946}},
{{8'sd-75, 13'sd-2289, 13'sd-2421}, {12'sd-1960, 12'sd1533, 12'sd-1538}, {13'sd-2195, 13'sd-2670, 13'sd-2548}},
{{13'sd-3251, 12'sd1254, 11'sd-678}, {12'sd2012, 12'sd-1577, 13'sd-2172}, {9'sd160, 12'sd1240, 13'sd-2486}},
{{11'sd-857, 13'sd-2510, 13'sd-2401}, {14'sd-4121, 12'sd-1959, 11'sd-940}, {13'sd-3979, 13'sd-2574, 11'sd-822}},
{{12'sd1255, 11'sd888, 11'sd901}, {12'sd-1698, 9'sd-174, 12'sd-1499}, {13'sd2431, 9'sd-135, 13'sd2733}},
{{7'sd-40, 13'sd-2956, 11'sd923}, {12'sd-1727, 13'sd-2915, 8'sd-123}, {13'sd-3569, 11'sd-790, 10'sd272}},
{{9'sd-204, 13'sd-2766, 13'sd2400}, {12'sd-1777, 12'sd-1368, 13'sd2194}, {12'sd1999, 12'sd2028, 9'sd-134}},
{{11'sd-699, 13'sd-2824, 13'sd-2818}, {11'sd-645, 11'sd-822, 12'sd-1771}, {13'sd-2288, 13'sd-2253, 12'sd-1105}},
{{13'sd-2395, 7'sd-50, 12'sd-1097}, {12'sd1615, 12'sd-1227, 12'sd-1740}, {12'sd1802, 13'sd2745, 11'sd777}},
{{11'sd777, 11'sd-824, 12'sd1773}, {13'sd-2145, 13'sd2438, 10'sd-453}, {10'sd-438, 12'sd-1672, 13'sd-2142}},
{{12'sd1626, 11'sd811, 6'sd-17}, {13'sd2283, 9'sd130, 12'sd-1592}, {9'sd134, 12'sd-1426, 5'sd-10}},
{{12'sd1880, 10'sd-470, 11'sd746}, {12'sd1141, 10'sd262, 10'sd-314}, {13'sd-2558, 13'sd-2272, 11'sd-670}},
{{12'sd1937, 8'sd70, 13'sd2710}, {11'sd552, 12'sd1887, 12'sd-1579}, {11'sd-736, 12'sd1339, 11'sd855}}},
{
{{13'sd-2373, 7'sd47, 12'sd-1333}, {12'sd-1190, 12'sd1314, 13'sd-2287}, {12'sd1996, 11'sd-936, 12'sd2042}},
{{11'sd599, 13'sd-2283, 11'sd907}, {11'sd929, 13'sd-2307, 11'sd-864}, {12'sd-2010, 11'sd645, 11'sd962}},
{{9'sd244, 12'sd-2016, 13'sd-2376}, {13'sd2127, 12'sd1432, 13'sd-2243}, {12'sd1510, 9'sd-149, 12'sd-1776}},
{{13'sd-2289, 12'sd1318, 13'sd2574}, {10'sd343, 13'sd2261, 11'sd815}, {12'sd-1797, 12'sd1179, 9'sd179}},
{{13'sd-2794, 13'sd-2184, 11'sd627}, {13'sd-2148, 13'sd-3743, 12'sd-1246}, {13'sd-3923, 12'sd-1369, 13'sd-3027}},
{{13'sd2205, 12'sd-1212, 11'sd649}, {13'sd2261, 11'sd-807, 12'sd-1208}, {12'sd-1766, 12'sd1144, 12'sd-1659}},
{{12'sd1563, 7'sd62, 11'sd-939}, {13'sd-2584, 13'sd-3170, 10'sd268}, {11'sd-645, 12'sd1431, 8'sd85}},
{{13'sd-2125, 13'sd-2490, 12'sd1647}, {10'sd348, 12'sd1301, 13'sd-2056}, {11'sd618, 12'sd-1333, 9'sd254}},
{{11'sd-962, 11'sd810, 13'sd2236}, {12'sd1748, 12'sd1906, 11'sd750}, {10'sd438, 12'sd1029, 13'sd-2387}},
{{11'sd-627, 13'sd-2147, 13'sd-3061}, {13'sd-2481, 13'sd2247, 12'sd-1765}, {9'sd223, 12'sd-1507, 11'sd-931}},
{{12'sd1891, 11'sd854, 12'sd-1030}, {13'sd-2826, 13'sd-3043, 12'sd1679}, {13'sd2466, 11'sd720, 13'sd-2673}},
{{12'sd1173, 12'sd2001, 12'sd1490}, {13'sd2293, 12'sd-1077, 13'sd2138}, {12'sd1885, 13'sd-2691, 12'sd-1116}},
{{11'sd-908, 13'sd-3082, 12'sd-1976}, {11'sd906, 13'sd-3553, 13'sd-2776}, {13'sd-2406, 11'sd648, 10'sd-496}},
{{11'sd-544, 13'sd2633, 13'sd2618}, {11'sd-969, 11'sd798, 11'sd819}, {12'sd1090, 13'sd2188, 13'sd-2624}},
{{12'sd1852, 12'sd1094, 7'sd37}, {12'sd1973, 10'sd322, 13'sd-2786}, {12'sd1268, 6'sd-16, 12'sd-1589}},
{{12'sd-1229, 12'sd-1802, 11'sd-877}, {12'sd1374, 11'sd782, 9'sd144}, {10'sd-367, 11'sd-701, 10'sd263}},
{{6'sd-16, 12'sd-1360, 12'sd1376}, {12'sd1536, 12'sd2005, 11'sd576}, {8'sd65, 7'sd-33, 11'sd-772}},
{{13'sd-2872, 13'sd-3369, 10'sd-504}, {11'sd-799, 13'sd-3019, 9'sd-218}, {13'sd-2748, 9'sd149, 8'sd-77}},
{{13'sd-2350, 11'sd541, 12'sd1884}, {12'sd-1290, 13'sd2130, 12'sd1275}, {12'sd1629, 13'sd-2253, 12'sd-1518}},
{{10'sd-274, 12'sd1714, 9'sd193}, {12'sd-1127, 10'sd296, 13'sd2395}, {13'sd2465, 13'sd-2087, 12'sd-1789}},
{{10'sd-323, 13'sd2848, 12'sd1071}, {11'sd-935, 12'sd-1709, 10'sd-324}, {11'sd-864, 12'sd-1062, 12'sd2008}},
{{11'sd-726, 10'sd-494, 9'sd238}, {13'sd-2183, 6'sd29, 10'sd-292}, {13'sd-2266, 12'sd-1648, 12'sd1111}},
{{10'sd328, 13'sd2441, 13'sd-2115}, {11'sd-842, 11'sd516, 9'sd244}, {12'sd-1157, 10'sd308, 11'sd-721}},
{{12'sd-1251, 9'sd183, 11'sd-557}, {11'sd524, 11'sd760, 12'sd-1393}, {13'sd-2293, 12'sd-1146, 13'sd2935}},
{{12'sd-1502, 11'sd-911, 12'sd1868}, {13'sd-2511, 12'sd1615, 12'sd1765}, {13'sd-2412, 11'sd776, 12'sd-1033}},
{{12'sd-1038, 12'sd1263, 12'sd-1614}, {13'sd-2440, 9'sd181, 11'sd-655}, {12'sd1770, 13'sd-3112, 11'sd883}},
{{11'sd-895, 3'sd-3, 12'sd-1495}, {11'sd-824, 13'sd-2894, 11'sd596}, {14'sd-4935, 13'sd-2076, 11'sd-581}},
{{11'sd760, 12'sd1715, 12'sd-1982}, {12'sd-1616, 13'sd2649, 11'sd-968}, {12'sd1621, 12'sd1587, 12'sd1858}},
{{10'sd-292, 13'sd-2164, 10'sd-421}, {13'sd2738, 11'sd-984, 10'sd-480}, {10'sd-463, 11'sd-945, 12'sd1841}},
{{5'sd12, 13'sd2118, 12'sd1363}, {10'sd-266, 11'sd-702, 11'sd-683}, {11'sd-575, 5'sd8, 12'sd1508}},
{{12'sd1967, 12'sd1189, 13'sd-2068}, {12'sd1646, 13'sd2546, 11'sd824}, {13'sd2065, 12'sd1750, 12'sd-1985}},
{{12'sd1402, 12'sd1148, 13'sd-2055}, {10'sd-448, 9'sd-249, 7'sd-36}, {12'sd-1647, 13'sd-2749, 11'sd-817}},
{{13'sd-2070, 12'sd-1624, 13'sd2209}, {12'sd1970, 12'sd-2031, 12'sd-1219}, {12'sd-1417, 11'sd-637, 10'sd-507}},
{{12'sd1883, 10'sd-305, 11'sd-733}, {12'sd-1404, 13'sd-2271, 12'sd-1837}, {12'sd1822, 11'sd774, 13'sd2384}},
{{13'sd-2580, 13'sd2495, 11'sd-764}, {13'sd2159, 13'sd3029, 10'sd278}, {12'sd-1403, 12'sd-1478, 12'sd-1496}},
{{10'sd366, 11'sd-948, 11'sd613}, {12'sd1425, 9'sd241, 12'sd1308}, {11'sd825, 13'sd2243, 12'sd1098}},
{{12'sd1495, 12'sd-1120, 12'sd1530}, {11'sd-739, 13'sd3576, 11'sd-902}, {10'sd-332, 13'sd2881, 13'sd2207}},
{{11'sd-930, 10'sd-488, 12'sd-1376}, {10'sd-488, 13'sd-3076, 13'sd-2729}, {13'sd2206, 12'sd-1655, 12'sd1802}},
{{12'sd-1496, 11'sd-606, 12'sd1146}, {13'sd-2599, 13'sd2505, 12'sd-1219}, {10'sd-385, 13'sd2357, 13'sd2286}},
{{13'sd2527, 12'sd-1458, 11'sd748}, {12'sd-1474, 13'sd2199, 11'sd836}, {11'sd-967, 13'sd-2574, 10'sd-379}},
{{10'sd313, 13'sd-2263, 11'sd-563}, {12'sd-2034, 12'sd1196, 13'sd-2988}, {11'sd612, 10'sd299, 13'sd2362}},
{{12'sd-1041, 11'sd805, 6'sd25}, {12'sd1309, 13'sd-3450, 13'sd-3407}, {10'sd466, 12'sd1303, 12'sd-1569}},
{{12'sd-1067, 12'sd1216, 10'sd454}, {12'sd1520, 13'sd2354, 2'sd1}, {12'sd-1855, 9'sd188, 13'sd2505}},
{{10'sd503, 13'sd-2542, 12'sd1869}, {13'sd-4065, 13'sd-3674, 12'sd-1969}, {14'sd-4119, 13'sd-2900, 13'sd-2860}},
{{12'sd1946, 13'sd2312, 13'sd-2638}, {12'sd-1518, 12'sd-1834, 12'sd1930}, {10'sd434, 7'sd-58, 10'sd-391}},
{{13'sd2496, 13'sd2849, 6'sd-21}, {12'sd-1478, 12'sd1474, 13'sd2197}, {12'sd1924, 9'sd150, 9'sd-245}},
{{12'sd1300, 12'sd1975, 13'sd-2207}, {10'sd292, 11'sd886, 12'sd1574}, {13'sd-2328, 12'sd-1466, 13'sd-2160}},
{{13'sd-2354, 12'sd-1849, 12'sd1168}, {12'sd1276, 11'sd902, 10'sd-265}, {11'sd-674, 10'sd390, 12'sd1610}},
{{4'sd7, 11'sd-699, 5'sd-9}, {11'sd-682, 13'sd2264, 13'sd2760}, {13'sd-2071, 13'sd3242, 13'sd3329}},
{{11'sd679, 13'sd3123, 9'sd203}, {13'sd3036, 12'sd1982, 9'sd185}, {12'sd1316, 13'sd3411, 12'sd1681}},
{{11'sd534, 13'sd2345, 13'sd2549}, {12'sd-1202, 8'sd-68, 12'sd1706}, {13'sd-2372, 12'sd-1409, 9'sd-238}},
{{12'sd-1714, 12'sd-1833, 9'sd-227}, {11'sd-544, 9'sd-152, 10'sd411}, {11'sd-873, 11'sd986, 6'sd27}},
{{11'sd922, 13'sd-2380, 13'sd2521}, {13'sd2667, 12'sd1433, 12'sd-1298}, {12'sd-1302, 10'sd-406, 12'sd1738}},
{{12'sd-1774, 11'sd-950, 13'sd-2555}, {12'sd-1617, 10'sd-343, 13'sd-2523}, {12'sd-1968, 12'sd-1660, 12'sd1048}},
{{13'sd-2338, 13'sd-2081, 12'sd-2037}, {13'sd-3293, 13'sd-3901, 12'sd-1766}, {13'sd-2525, 11'sd688, 12'sd-1864}},
{{12'sd-2004, 11'sd640, 11'sd-540}, {10'sd-362, 10'sd335, 12'sd-1736}, {13'sd2709, 13'sd3177, 11'sd736}},
{{13'sd-2181, 13'sd-2268, 14'sd-4345}, {8'sd95, 11'sd990, 13'sd-4072}, {13'sd-3162, 13'sd-2442, 10'sd405}},
{{12'sd1351, 11'sd767, 12'sd-1107}, {10'sd358, 12'sd1431, 13'sd-2796}, {12'sd-1170, 12'sd1867, 13'sd-2818}},
{{12'sd-1103, 12'sd-1478, 11'sd-646}, {13'sd-2632, 8'sd124, 13'sd-2135}, {9'sd-145, 10'sd374, 13'sd-2876}},
{{11'sd530, 6'sd-23, 10'sd-326}, {12'sd1471, 12'sd1484, 11'sd-693}, {12'sd1316, 13'sd2518, 12'sd-2015}},
{{13'sd2425, 12'sd-1234, 10'sd-258}, {12'sd1581, 12'sd2032, 11'sd607}, {13'sd2434, 12'sd1135, 11'sd924}},
{{12'sd-1731, 12'sd-1216, 11'sd939}, {10'sd-284, 10'sd-375, 11'sd608}, {12'sd1602, 10'sd-387, 11'sd-608}},
{{11'sd781, 13'sd2780, 12'sd1139}, {9'sd171, 11'sd-1001, 12'sd-1130}, {13'sd-3135, 9'sd198, 12'sd-1884}},
{{13'sd2801, 13'sd2351, 12'sd1042}, {12'sd1888, 10'sd488, 13'sd3182}, {13'sd3668, 12'sd1364, 12'sd1934}}},
{
{{12'sd1610, 9'sd-142, 10'sd326}, {10'sd-261, 10'sd-406, 11'sd842}, {13'sd2437, 12'sd1100, 12'sd-1143}},
{{13'sd-2144, 11'sd787, 10'sd-434}, {12'sd-1395, 12'sd2023, 12'sd-1494}, {9'sd-246, 11'sd-856, 12'sd-1326}},
{{11'sd-625, 11'sd-549, 13'sd2772}, {12'sd-1461, 13'sd2179, 11'sd515}, {12'sd1093, 13'sd2645, 13'sd2286}},
{{13'sd-2652, 13'sd-2682, 9'sd-228}, {13'sd-2731, 11'sd710, 12'sd-1767}, {12'sd1816, 11'sd544, 11'sd-759}},
{{13'sd2208, 7'sd45, 12'sd1762}, {13'sd-2931, 12'sd-1157, 12'sd1523}, {13'sd-2550, 9'sd-169, 13'sd-2959}},
{{11'sd636, 12'sd1248, 13'sd3464}, {12'sd-1644, 12'sd1881, 12'sd-1409}, {13'sd2084, 11'sd796, 12'sd-1678}},
{{13'sd-3368, 11'sd678, 9'sd180}, {10'sd293, 10'sd460, 13'sd-2105}, {11'sd723, 12'sd-1373, 12'sd1209}},
{{11'sd-919, 12'sd1128, 12'sd-1578}, {9'sd-243, 11'sd917, 13'sd2352}, {12'sd-2030, 10'sd442, 10'sd508}},
{{12'sd1733, 11'sd-579, 13'sd2150}, {12'sd1834, 12'sd-1988, 12'sd-1993}, {13'sd-2377, 13'sd-2911, 7'sd-59}},
{{13'sd2105, 12'sd1555, 4'sd-6}, {12'sd-1561, 12'sd-1672, 11'sd-888}, {11'sd-734, 12'sd-1507, 13'sd2095}},
{{11'sd719, 11'sd-603, 10'sd-458}, {12'sd1376, 11'sd-737, 13'sd-2204}, {10'sd-399, 12'sd1070, 10'sd-274}},
{{13'sd2111, 13'sd-2108, 11'sd890}, {12'sd1331, 12'sd-1557, 13'sd2597}, {13'sd-2566, 11'sd907, 11'sd-858}},
{{10'sd-384, 13'sd2199, 13'sd-3051}, {12'sd1267, 13'sd-2863, 11'sd-715}, {13'sd2201, 12'sd1459, 3'sd3}},
{{13'sd2064, 11'sd-647, 12'sd1385}, {12'sd1207, 11'sd714, 13'sd-2555}, {9'sd169, 1'sd0, 11'sd591}},
{{9'sd238, 7'sd-45, 12'sd-1929}, {11'sd-804, 6'sd27, 12'sd1591}, {12'sd1890, 9'sd-184, 11'sd-1022}},
{{12'sd1284, 13'sd-2638, 11'sd671}, {13'sd2226, 13'sd2225, 12'sd1746}, {11'sd-567, 12'sd1539, 12'sd-1852}},
{{13'sd2340, 13'sd2530, 9'sd252}, {12'sd1499, 11'sd-780, 12'sd-1978}, {8'sd-103, 11'sd-805, 12'sd-1503}},
{{12'sd-1522, 12'sd1874, 10'sd332}, {12'sd-1629, 12'sd1863, 13'sd-2955}, {5'sd13, 12'sd-2029, 12'sd-1567}},
{{9'sd155, 10'sd-355, 12'sd1309}, {12'sd-1553, 13'sd2409, 13'sd2216}, {13'sd2223, 11'sd-573, 13'sd2344}},
{{12'sd-1952, 11'sd913, 13'sd2221}, {13'sd2561, 12'sd1201, 11'sd609}, {13'sd-2654, 13'sd2347, 12'sd1603}},
{{12'sd-1312, 11'sd636, 13'sd2320}, {10'sd-285, 9'sd-184, 13'sd2280}, {11'sd1007, 12'sd-1214, 12'sd1275}},
{{9'sd133, 12'sd-1979, 9'sd204}, {7'sd-38, 12'sd-2038, 8'sd68}, {12'sd2007, 12'sd1074, 12'sd-1829}},
{{12'sd1462, 10'sd-494, 13'sd2204}, {10'sd483, 12'sd1304, 12'sd-1691}, {6'sd-30, 12'sd1482, 12'sd-1993}},
{{12'sd1639, 12'sd1508, 13'sd2227}, {13'sd-2170, 12'sd1866, 11'sd-863}, {10'sd-463, 7'sd41, 6'sd19}},
{{11'sd-605, 12'sd1497, 13'sd2087}, {12'sd-1821, 13'sd-2492, 12'sd-1278}, {13'sd-2478, 11'sd680, 11'sd-974}},
{{13'sd2717, 9'sd-182, 11'sd-1015}, {12'sd1067, 12'sd-1404, 12'sd1395}, {9'sd178, 12'sd1468, 12'sd1633}},
{{9'sd242, 10'sd371, 11'sd819}, {13'sd-2613, 11'sd877, 12'sd-1926}, {10'sd-465, 11'sd543, 10'sd322}},
{{12'sd1959, 12'sd-1359, 11'sd-966}, {11'sd-791, 12'sd-1304, 12'sd-1102}, {12'sd-1297, 10'sd371, 12'sd-1584}},
{{12'sd1808, 12'sd-1923, 10'sd-505}, {13'sd2714, 12'sd1422, 12'sd-1434}, {11'sd678, 12'sd-1698, 12'sd1718}},
{{12'sd1346, 13'sd2177, 12'sd-1342}, {8'sd123, 11'sd-642, 9'sd243}, {9'sd-171, 13'sd-2403, 13'sd3007}},
{{10'sd-321, 12'sd1319, 11'sd895}, {9'sd-152, 12'sd-1166, 12'sd1560}, {12'sd-1535, 13'sd-2503, 9'sd-227}},
{{11'sd-662, 12'sd-1791, 13'sd-2614}, {13'sd2528, 9'sd-131, 12'sd1182}, {12'sd1685, 12'sd1986, 12'sd-1433}},
{{12'sd-1384, 12'sd1669, 11'sd-727}, {9'sd134, 12'sd-1282, 12'sd-1401}, {13'sd-2977, 11'sd-686, 10'sd377}},
{{12'sd-1700, 13'sd2877, 13'sd2329}, {11'sd-697, 12'sd-1885, 8'sd-94}, {12'sd1113, 12'sd1501, 12'sd1668}},
{{9'sd-230, 12'sd-1037, 11'sd558}, {12'sd1539, 12'sd-1146, 13'sd2394}, {11'sd658, 11'sd757, 13'sd2718}},
{{13'sd-2262, 12'sd1308, 13'sd2202}, {12'sd1302, 11'sd-630, 9'sd-134}, {12'sd1548, 13'sd2049, 13'sd2136}},
{{10'sd428, 12'sd1890, 13'sd2055}, {11'sd612, 13'sd3099, 7'sd-41}, {13'sd-2168, 12'sd-1466, 9'sd215}},
{{11'sd607, 12'sd1870, 11'sd-601}, {10'sd403, 10'sd-287, 13'sd-2078}, {8'sd93, 12'sd-1721, 13'sd-3025}},
{{12'sd1331, 11'sd947, 13'sd2109}, {11'sd-543, 11'sd-846, 13'sd-2249}, {11'sd-618, 11'sd643, 11'sd643}},
{{11'sd-583, 12'sd-1684, 13'sd-2479}, {12'sd1340, 10'sd-328, 13'sd-2638}, {13'sd2320, 11'sd-671, 12'sd-1236}},
{{12'sd1152, 12'sd-1951, 7'sd-33}, {12'sd1954, 11'sd773, 13'sd2220}, {13'sd-2891, 10'sd-319, 12'sd-1962}},
{{12'sd-1029, 12'sd-1213, 13'sd-2105}, {11'sd872, 10'sd-322, 12'sd-1741}, {12'sd1576, 12'sd1405, 11'sd-648}},
{{11'sd894, 12'sd1050, 13'sd2239}, {13'sd2887, 11'sd-560, 13'sd2174}, {12'sd-1450, 9'sd155, 11'sd-837}},
{{12'sd-1905, 13'sd-2175, 12'sd-2015}, {13'sd-3372, 11'sd-969, 13'sd-2407}, {13'sd-3054, 12'sd-1206, 13'sd2237}},
{{12'sd-1916, 13'sd2235, 12'sd1091}, {11'sd-855, 11'sd620, 12'sd1667}, {10'sd335, 13'sd-2639, 12'sd1342}},
{{12'sd1997, 13'sd2568, 12'sd-1675}, {12'sd-1198, 12'sd1613, 12'sd-1151}, {12'sd1506, 10'sd-461, 12'sd-1158}},
{{12'sd1923, 13'sd2235, 12'sd1272}, {11'sd694, 13'sd-2268, 9'sd-231}, {13'sd-2286, 13'sd2798, 12'sd1267}},
{{9'sd132, 10'sd-397, 13'sd-2557}, {12'sd-1538, 12'sd-2031, 12'sd-1395}, {12'sd1282, 12'sd-1858, 12'sd2013}},
{{7'sd53, 8'sd-78, 11'sd-573}, {12'sd1160, 11'sd-775, 11'sd-661}, {13'sd2953, 11'sd669, 13'sd2612}},
{{12'sd-1958, 12'sd1583, 13'sd2757}, {12'sd-1084, 11'sd525, 11'sd909}, {13'sd2096, 10'sd262, 11'sd610}},
{{11'sd707, 12'sd1301, 12'sd-1194}, {10'sd-313, 12'sd-1836, 11'sd740}, {13'sd-2593, 12'sd1840, 13'sd-2360}},
{{12'sd1621, 12'sd-1687, 11'sd-883}, {11'sd541, 13'sd-2455, 13'sd-2302}, {12'sd1338, 13'sd-2355, 9'sd248}},
{{13'sd2816, 12'sd-1442, 13'sd-2242}, {12'sd-1317, 11'sd664, 6'sd-23}, {12'sd1325, 11'sd-739, 11'sd587}},
{{11'sd-555, 12'sd1525, 12'sd1962}, {13'sd-2510, 12'sd1160, 12'sd1487}, {8'sd99, 12'sd-1104, 12'sd1322}},
{{13'sd-2717, 12'sd-1643, 12'sd-1554}, {13'sd-2200, 13'sd-2194, 11'sd676}, {12'sd-1405, 10'sd-275, 12'sd-1478}},
{{11'sd-747, 13'sd2280, 13'sd2755}, {11'sd-517, 11'sd761, 13'sd2146}, {13'sd2355, 12'sd-1116, 11'sd-825}},
{{10'sd-423, 8'sd118, 13'sd-2986}, {9'sd221, 8'sd-94, 13'sd-3295}, {8'sd-100, 12'sd-1930, 13'sd-2864}},
{{9'sd-133, 12'sd1593, 12'sd-1275}, {8'sd-90, 12'sd1706, 13'sd-2095}, {10'sd374, 10'sd-432, 12'sd-1683}},
{{11'sd-1004, 13'sd2446, 11'sd-864}, {12'sd1738, 11'sd950, 12'sd-1190}, {13'sd-2337, 13'sd-2420, 11'sd871}},
{{12'sd1053, 12'sd-1444, 12'sd-1485}, {12'sd1050, 12'sd1914, 12'sd1530}, {11'sd748, 13'sd2667, 7'sd-49}},
{{11'sd-517, 12'sd1049, 13'sd2079}, {12'sd-1444, 12'sd-1446, 13'sd-2693}, {9'sd240, 11'sd804, 12'sd1289}},
{{12'sd1652, 12'sd1529, 9'sd-154}, {11'sd-693, 12'sd-1357, 10'sd-267}, {11'sd-964, 8'sd75, 5'sd-9}},
{{10'sd309, 13'sd2308, 12'sd-1090}, {11'sd-722, 12'sd-1823, 13'sd-2280}, {13'sd-2276, 12'sd-1508, 12'sd1275}},
{{11'sd-617, 10'sd368, 13'sd-2372}, {6'sd-23, 13'sd2140, 12'sd-1510}, {11'sd894, 12'sd-1434, 11'sd633}}},
{
{{11'sd993, 13'sd2332, 11'sd-951}, {12'sd1983, 12'sd1026, 13'sd-2437}, {12'sd-1111, 9'sd-249, 13'sd2240}},
{{11'sd-829, 10'sd511, 13'sd-2109}, {9'sd-193, 11'sd565, 10'sd-313}, {10'sd-376, 12'sd1868, 12'sd-1669}},
{{8'sd106, 11'sd-1000, 13'sd3265}, {6'sd24, 13'sd-2590, 12'sd-1604}, {13'sd-2236, 13'sd2304, 13'sd2378}},
{{12'sd-1341, 12'sd-1889, 13'sd-2508}, {12'sd1662, 12'sd-1816, 13'sd2056}, {13'sd-2407, 11'sd696, 12'sd1299}},
{{13'sd3360, 12'sd1478, 14'sd4933}, {14'sd4909, 14'sd5233, 9'sd157}, {12'sd1611, 8'sd75, 9'sd-135}},
{{12'sd1384, 11'sd-932, 10'sd-342}, {11'sd829, 12'sd-1439, 11'sd540}, {10'sd-476, 11'sd-728, 11'sd596}},
{{13'sd2780, 10'sd-346, 13'sd2492}, {12'sd1160, 12'sd-1147, 13'sd-2083}, {12'sd-1323, 10'sd-498, 14'sd-4333}},
{{11'sd649, 12'sd-1177, 13'sd-2630}, {8'sd82, 12'sd-1122, 13'sd2140}, {8'sd-70, 12'sd-1761, 11'sd-981}},
{{11'sd932, 12'sd-1253, 12'sd-1578}, {13'sd-2070, 12'sd-1931, 13'sd2459}, {10'sd-476, 12'sd-1025, 12'sd-1736}},
{{8'sd108, 12'sd-1768, 12'sd-1759}, {11'sd777, 12'sd-1694, 12'sd1556}, {11'sd905, 9'sd197, 11'sd724}},
{{13'sd2462, 13'sd2964, 10'sd429}, {13'sd-2817, 4'sd-7, 12'sd1140}, {8'sd106, 13'sd-2606, 11'sd-681}},
{{12'sd1876, 13'sd2770, 13'sd2603}, {13'sd2622, 11'sd672, 13'sd2405}, {11'sd-971, 7'sd-34, 13'sd2662}},
{{13'sd-3531, 9'sd-237, 12'sd-1713}, {12'sd-1340, 13'sd-2323, 9'sd196}, {14'sd-4457, 12'sd-1309, 12'sd1328}},
{{11'sd593, 12'sd1909, 13'sd-2799}, {12'sd-1923, 6'sd22, 11'sd-554}, {11'sd-603, 11'sd-747, 12'sd1332}},
{{14'sd4431, 14'sd5585, 14'sd4906}, {13'sd2439, 13'sd3495, 13'sd3376}, {14'sd7305, 12'sd-1444, 12'sd-1367}},
{{13'sd-3445, 11'sd-894, 13'sd-2776}, {12'sd1742, 12'sd1104, 13'sd-2067}, {12'sd1119, 11'sd-618, 13'sd-3148}},
{{13'sd-2982, 11'sd-800, 13'sd-3256}, {11'sd-966, 13'sd2646, 10'sd321}, {12'sd-1233, 11'sd698, 11'sd-663}},
{{7'sd-33, 12'sd1462, 13'sd2538}, {10'sd-422, 11'sd-631, 12'sd1088}, {7'sd-54, 12'sd-1755, 11'sd-526}},
{{13'sd2345, 10'sd300, 13'sd-3032}, {11'sd-728, 11'sd615, 12'sd1885}, {12'sd1967, 12'sd1569, 13'sd-2959}},
{{12'sd1036, 12'sd1670, 10'sd-366}, {11'sd744, 10'sd465, 11'sd600}, {12'sd1137, 12'sd-1689, 12'sd1275}},
{{13'sd3311, 11'sd579, 12'sd1079}, {9'sd206, 12'sd-1524, 8'sd85}, {11'sd-849, 12'sd1440, 11'sd-927}},
{{12'sd-1411, 10'sd454, 11'sd-893}, {12'sd-1079, 12'sd-1149, 12'sd1147}, {12'sd1034, 12'sd-1245, 13'sd2147}},
{{13'sd-2670, 13'sd2189, 13'sd-2709}, {12'sd-1630, 12'sd1160, 11'sd-793}, {10'sd-491, 12'sd1843, 12'sd-1664}},
{{12'sd1052, 12'sd-1976, 11'sd863}, {13'sd2451, 13'sd-2543, 10'sd-505}, {9'sd153, 9'sd162, 11'sd737}},
{{9'sd-214, 11'sd-793, 13'sd-2462}, {13'sd2232, 13'sd-2505, 13'sd-2566}, {13'sd-3008, 13'sd-3052, 12'sd-2040}},
{{12'sd-1033, 12'sd1452, 13'sd2561}, {12'sd-1881, 11'sd-785, 11'sd-715}, {8'sd-120, 13'sd-2817, 12'sd-1723}},
{{13'sd-2444, 14'sd-4164, 13'sd-2773}, {13'sd-2675, 14'sd-5238, 12'sd1412}, {14'sd-6871, 14'sd-4525, 10'sd257}},
{{12'sd1444, 13'sd2197, 10'sd-458}, {12'sd1290, 12'sd1140, 13'sd2892}, {12'sd1528, 13'sd-2145, 12'sd-1803}},
{{7'sd-53, 11'sd-806, 11'sd-567}, {12'sd-1609, 12'sd1105, 13'sd-2409}, {13'sd-4065, 12'sd-1376, 9'sd-174}},
{{11'sd-522, 11'sd-926, 13'sd2582}, {12'sd1063, 12'sd1564, 11'sd-670}, {13'sd-2601, 12'sd-1759, 13'sd3012}},
{{8'sd79, 12'sd-1678, 13'sd-2481}, {12'sd1849, 13'sd-2064, 12'sd-1260}, {13'sd2773, 10'sd-307, 12'sd1199}},
{{10'sd258, 13'sd2607, 12'sd1857}, {12'sd-1689, 13'sd2177, 8'sd-126}, {12'sd-1954, 11'sd-977, 11'sd-895}},
{{11'sd-942, 12'sd1598, 12'sd1802}, {9'sd-205, 11'sd611, 9'sd-144}, {8'sd68, 12'sd1504, 10'sd314}},
{{13'sd2991, 12'sd1872, 12'sd-1520}, {11'sd582, 12'sd1741, 13'sd-2403}, {13'sd2753, 12'sd1483, 8'sd102}},
{{5'sd-12, 11'sd-547, 13'sd-2542}, {9'sd-238, 13'sd2171, 11'sd-750}, {12'sd-1220, 13'sd2909, 9'sd-164}},
{{10'sd-433, 12'sd1871, 11'sd828}, {12'sd-1690, 12'sd-1095, 12'sd-1049}, {12'sd-1088, 12'sd1068, 13'sd-2781}},
{{14'sd-4660, 13'sd-3163, 14'sd-4685}, {13'sd-3100, 11'sd-1004, 11'sd-931}, {13'sd-3611, 10'sd-320, 11'sd-627}},
{{12'sd1461, 13'sd2752, 13'sd2252}, {12'sd-1331, 9'sd194, 13'sd2321}, {12'sd-1460, 12'sd-1952, 5'sd13}},
{{10'sd441, 12'sd-1910, 10'sd-265}, {8'sd118, 13'sd-2071, 12'sd1782}, {13'sd2338, 9'sd-186, 9'sd250}},
{{12'sd1419, 10'sd267, 11'sd-540}, {13'sd-2128, 11'sd-817, 9'sd-230}, {11'sd907, 13'sd2290, 12'sd1029}},
{{13'sd2294, 8'sd90, 13'sd3040}, {10'sd391, 11'sd1023, 12'sd-1886}, {13'sd-2195, 8'sd-74, 12'sd-1871}},
{{12'sd2012, 11'sd966, 11'sd668}, {12'sd1906, 11'sd-1001, 12'sd1805}, {10'sd418, 12'sd1429, 13'sd2511}},
{{13'sd-2063, 12'sd-1074, 10'sd-349}, {13'sd-3468, 13'sd-2263, 11'sd968}, {12'sd-1073, 12'sd1773, 12'sd-1648}},
{{13'sd-2761, 12'sd1647, 8'sd-114}, {13'sd-4095, 12'sd1033, 11'sd686}, {15'sd-8522, 10'sd435, 11'sd613}},
{{12'sd-1259, 12'sd-1163, 8'sd-70}, {11'sd-782, 13'sd-2757, 12'sd-1912}, {9'sd177, 12'sd-1999, 12'sd-2040}},
{{12'sd1176, 8'sd119, 13'sd-2238}, {11'sd983, 12'sd-1110, 13'sd2240}, {13'sd2838, 12'sd2008, 12'sd-1656}},
{{13'sd-3322, 13'sd-3808, 12'sd-1690}, {11'sd892, 12'sd-1637, 12'sd1609}, {10'sd260, 11'sd-665, 11'sd581}},
{{12'sd1078, 10'sd390, 12'sd2022}, {12'sd-1076, 11'sd812, 11'sd728}, {13'sd2164, 9'sd-154, 12'sd1184}},
{{12'sd-1395, 12'sd-1588, 13'sd2163}, {11'sd-994, 12'sd-1691, 13'sd2630}, {10'sd479, 12'sd-1786, 10'sd-327}},
{{12'sd1824, 8'sd79, 11'sd-935}, {13'sd2464, 11'sd632, 13'sd-2360}, {12'sd1309, 11'sd-988, 10'sd402}},
{{13'sd2061, 12'sd-1605, 11'sd-672}, {10'sd504, 13'sd2220, 12'sd1469}, {13'sd2136, 12'sd-1822, 10'sd351}},
{{13'sd2390, 12'sd-1153, 11'sd-779}, {13'sd-2349, 12'sd1522, 10'sd-464}, {12'sd-1554, 13'sd2142, 11'sd-867}},
{{13'sd3029, 13'sd3368, 13'sd3784}, {11'sd-625, 2'sd-1, 13'sd2584}, {12'sd1922, 13'sd3180, 13'sd-2685}},
{{13'sd-2472, 13'sd-2699, 12'sd1930}, {7'sd-57, 13'sd-2380, 13'sd-3013}, {12'sd-1655, 12'sd-1682, 13'sd-2700}},
{{11'sd716, 12'sd1482, 11'sd-680}, {12'sd1536, 13'sd-2659, 12'sd1756}, {13'sd2068, 13'sd-2649, 10'sd264}},
{{13'sd-2596, 13'sd-3101, 11'sd618}, {11'sd-535, 13'sd2215, 11'sd-717}, {10'sd303, 13'sd2584, 12'sd1545}},
{{13'sd2919, 12'sd-1742, 12'sd1404}, {9'sd-175, 11'sd-872, 11'sd-659}, {14'sd7078, 13'sd2535, 10'sd353}},
{{11'sd-861, 12'sd-1724, 13'sd2436}, {11'sd-645, 11'sd-518, 10'sd-371}, {11'sd-636, 12'sd1266, 12'sd-1891}},
{{10'sd506, 11'sd715, 12'sd-1243}, {10'sd-453, 13'sd2607, 11'sd-625}, {12'sd1033, 12'sd1703, 10'sd262}},
{{11'sd543, 11'sd931, 13'sd2338}, {12'sd-1563, 13'sd3069, 11'sd-818}, {12'sd-1359, 12'sd-1308, 9'sd246}},
{{13'sd-2228, 10'sd419, 12'sd-1566}, {12'sd2020, 13'sd2382, 12'sd-1228}, {8'sd92, 11'sd-752, 8'sd110}},
{{7'sd38, 10'sd436, 13'sd-2642}, {11'sd-848, 11'sd750, 11'sd838}, {8'sd89, 11'sd-625, 12'sd-1550}},
{{12'sd1880, 7'sd57, 12'sd-1795}, {12'sd1720, 10'sd349, 13'sd2171}, {10'sd381, 12'sd1212, 11'sd566}},
{{13'sd2257, 12'sd-1187, 13'sd3301}, {11'sd806, 11'sd774, 8'sd73}, {12'sd-1780, 9'sd-175, 12'sd-1314}}},
{
{{12'sd-1125, 10'sd-320, 13'sd-2296}, {12'sd1830, 12'sd1951, 12'sd-1178}, {11'sd939, 12'sd1553, 10'sd-338}},
{{13'sd2299, 10'sd257, 12'sd1715}, {11'sd1014, 12'sd-1906, 13'sd-3869}, {13'sd-2848, 11'sd604, 13'sd-3007}},
{{5'sd-10, 13'sd-2239, 12'sd1652}, {13'sd-3018, 12'sd1881, 12'sd1551}, {13'sd-3784, 11'sd827, 11'sd734}},
{{13'sd2078, 12'sd-1247, 11'sd585}, {13'sd2625, 13'sd2887, 12'sd-1252}, {13'sd-2477, 12'sd1234, 12'sd1178}},
{{12'sd1298, 11'sd535, 12'sd-1626}, {13'sd2455, 14'sd4352, 11'sd841}, {13'sd2053, 9'sd205, 13'sd2356}},
{{11'sd817, 13'sd2823, 11'sd543}, {11'sd-709, 12'sd1302, 14'sd5239}, {11'sd759, 14'sd4626, 14'sd4960}},
{{14'sd7197, 13'sd2703, 13'sd3800}, {14'sd4117, 14'sd6283, 13'sd3287}, {13'sd-3286, 13'sd-2162, 9'sd243}},
{{13'sd3074, 13'sd-2240, 11'sd-952}, {12'sd1182, 13'sd2306, 13'sd-2104}, {8'sd-81, 13'sd2400, 11'sd-548}},
{{12'sd1501, 13'sd-2613, 12'sd1671}, {12'sd1641, 12'sd-1796, 12'sd-1256}, {6'sd29, 9'sd-183, 13'sd-2817}},
{{12'sd-1217, 4'sd7, 13'sd2734}, {12'sd1417, 11'sd534, 11'sd-727}, {12'sd1417, 10'sd261, 11'sd-714}},
{{11'sd-707, 12'sd-1724, 13'sd2876}, {11'sd-551, 7'sd-55, 13'sd3893}, {14'sd-4535, 13'sd-4009, 11'sd-790}},
{{9'sd242, 9'sd211, 13'sd-2796}, {7'sd55, 13'sd-2404, 12'sd1474}, {10'sd-501, 12'sd-1170, 13'sd-2127}},
{{12'sd-1785, 12'sd1641, 11'sd688}, {9'sd154, 12'sd-1322, 9'sd-250}, {13'sd-2569, 13'sd-3337, 12'sd1337}},
{{11'sd-782, 12'sd-1299, 10'sd324}, {11'sd-906, 12'sd-1049, 11'sd-595}, {11'sd592, 11'sd639, 8'sd-87}},
{{11'sd-836, 13'sd3485, 13'sd3999}, {14'sd-5786, 12'sd1449, 13'sd2927}, {13'sd4042, 14'sd4930, 15'sd9164}},
{{12'sd-1300, 12'sd1086, 11'sd-952}, {13'sd2362, 12'sd1247, 6'sd23}, {13'sd-2376, 12'sd1227, 9'sd217}},
{{12'sd-1754, 13'sd-2248, 12'sd-1372}, {8'sd-99, 12'sd-1366, 12'sd-1244}, {11'sd799, 9'sd-188, 12'sd1486}},
{{9'sd134, 12'sd1983, 9'sd-205}, {13'sd-2439, 11'sd618, 12'sd1039}, {11'sd983, 11'sd-535, 13'sd2074}},
{{12'sd1399, 12'sd1581, 10'sd-474}, {11'sd-721, 13'sd-3109, 12'sd-1096}, {12'sd-1533, 12'sd-1966, 12'sd1810}},
{{12'sd1278, 12'sd1208, 10'sd296}, {13'sd2558, 13'sd2200, 13'sd-2425}, {12'sd1728, 12'sd-1191, 11'sd-811}},
{{11'sd514, 12'sd1426, 10'sd273}, {13'sd2535, 12'sd-1434, 11'sd929}, {13'sd2296, 13'sd2225, 11'sd549}},
{{13'sd2694, 10'sd503, 12'sd-1148}, {13'sd2260, 12'sd1929, 12'sd1138}, {7'sd-58, 11'sd531, 12'sd1165}},
{{11'sd841, 13'sd-3125, 11'sd-840}, {12'sd-1726, 13'sd-2574, 13'sd-3791}, {12'sd-2016, 13'sd2193, 11'sd-524}},
{{9'sd-236, 12'sd-1634, 11'sd-622}, {12'sd-1336, 12'sd1147, 13'sd-3162}, {12'sd-1131, 13'sd-3783, 12'sd-1556}},
{{11'sd827, 13'sd-2608, 7'sd32}, {12'sd-1691, 13'sd-2941, 12'sd-1665}, {11'sd-560, 12'sd1157, 13'sd2175}},
{{8'sd107, 12'sd-1077, 12'sd-1171}, {10'sd-424, 12'sd-1832, 13'sd2480}, {13'sd-2696, 9'sd-215, 11'sd638}},
{{10'sd-474, 13'sd-2363, 11'sd904}, {14'sd-4725, 14'sd-4884, 13'sd-3166}, {13'sd-3877, 14'sd-7130, 14'sd-5875}},
{{12'sd-1414, 11'sd617, 10'sd396}, {12'sd1060, 13'sd2334, 13'sd2818}, {13'sd2508, 12'sd1547, 13'sd3495}},
{{10'sd335, 12'sd-1400, 13'sd3082}, {14'sd-4141, 11'sd550, 12'sd1258}, {13'sd-4005, 13'sd-3764, 12'sd1775}},
{{12'sd-1627, 12'sd1902, 11'sd-767}, {12'sd1968, 13'sd-2605, 12'sd-2005}, {13'sd-3399, 11'sd-783, 14'sd-4785}},
{{13'sd2687, 13'sd-2594, 10'sd310}, {9'sd-214, 12'sd-1635, 11'sd-768}, {11'sd-625, 12'sd-1758, 12'sd1527}},
{{12'sd-1782, 13'sd2245, 9'sd-237}, {12'sd1288, 13'sd3399, 12'sd-1535}, {13'sd2186, 12'sd-1467, 13'sd3039}},
{{12'sd-2023, 11'sd817, 12'sd1423}, {13'sd-2296, 12'sd-1783, 13'sd2541}, {11'sd1019, 11'sd-620, 11'sd555}},
{{12'sd-1958, 13'sd-2242, 12'sd-1411}, {13'sd-2798, 10'sd357, 10'sd369}, {13'sd3087, 11'sd867, 9'sd142}},
{{12'sd1283, 11'sd868, 13'sd-3142}, {12'sd1241, 12'sd-2037, 12'sd-1505}, {12'sd1105, 13'sd2496, 14'sd-5073}},
{{11'sd851, 10'sd-503, 13'sd-2348}, {12'sd1313, 12'sd-1511, 12'sd2004}, {12'sd1463, 12'sd1699, 12'sd1103}},
{{13'sd3423, 10'sd-479, 12'sd-1354}, {13'sd2576, 13'sd3522, 11'sd728}, {11'sd-991, 14'sd4527, 12'sd1508}},
{{12'sd1264, 12'sd-1436, 13'sd3040}, {11'sd-968, 13'sd2675, 11'sd-797}, {12'sd1672, 10'sd405, 12'sd-1187}},
{{12'sd1774, 9'sd203, 13'sd2129}, {12'sd-1645, 11'sd883, 12'sd1893}, {12'sd-1214, 12'sd-1618, 13'sd-3415}},
{{12'sd1506, 12'sd-1841, 10'sd-491}, {12'sd1691, 12'sd-1990, 11'sd949}, {13'sd-2194, 12'sd1470, 13'sd2484}},
{{14'sd5584, 13'sd2419, 14'sd4224}, {9'sd185, 10'sd-265, 10'sd272}, {12'sd1532, 13'sd3246, 13'sd3845}},
{{12'sd-1032, 13'sd-2795, 10'sd489}, {8'sd77, 10'sd-484, 13'sd2125}, {11'sd-972, 11'sd-1010, 14'sd-4874}},
{{12'sd-1611, 11'sd748, 10'sd-379}, {12'sd-1543, 11'sd-766, 14'sd4180}, {13'sd-4065, 14'sd-5100, 10'sd-507}},
{{13'sd3602, 13'sd2142, 13'sd-2436}, {13'sd2766, 7'sd-35, 9'sd135}, {14'sd-6764, 12'sd-1300, 14'sd-7445}},
{{9'sd202, 13'sd2902, 12'sd1344}, {8'sd-115, 10'sd268, 13'sd-2810}, {12'sd1178, 10'sd319, 13'sd-2610}},
{{9'sd-249, 10'sd-362, 11'sd-876}, {9'sd-179, 11'sd598, 12'sd1167}, {12'sd-1576, 12'sd-1467, 11'sd594}},
{{11'sd-654, 13'sd-2413, 13'sd-2202}, {13'sd-4079, 12'sd-1135, 13'sd-3059}, {10'sd423, 12'sd1628, 13'sd-3055}},
{{12'sd-1659, 12'sd-1319, 8'sd-71}, {12'sd-1346, 11'sd934, 11'sd-660}, {11'sd986, 13'sd-2250, 13'sd-2438}},
{{13'sd-2412, 12'sd1204, 13'sd2940}, {12'sd-1399, 12'sd1714, 12'sd1692}, {9'sd232, 11'sd-667, 11'sd795}},
{{12'sd1367, 8'sd-100, 12'sd1272}, {13'sd-2581, 8'sd108, 13'sd-3387}, {13'sd2557, 10'sd-331, 11'sd-527}},
{{10'sd312, 12'sd1093, 12'sd1850}, {13'sd-2423, 12'sd-1226, 12'sd-1313}, {12'sd1864, 12'sd-1099, 11'sd885}},
{{12'sd1991, 13'sd-2379, 12'sd-1648}, {12'sd1600, 7'sd-63, 13'sd2918}, {11'sd-826, 12'sd1972, 5'sd-13}},
{{12'sd-1556, 10'sd-354, 8'sd121}, {11'sd1008, 14'sd5274, 13'sd3914}, {10'sd467, 10'sd-438, 11'sd995}},
{{12'sd1061, 12'sd1525, 13'sd-3121}, {12'sd1289, 12'sd-1045, 13'sd-2230}, {12'sd-1904, 12'sd-1783, 10'sd-401}},
{{13'sd-2721, 12'sd1752, 13'sd2929}, {12'sd-1568, 12'sd1175, 13'sd2854}, {13'sd-2599, 13'sd-3065, 11'sd-851}},
{{13'sd3291, 13'sd2295, 12'sd-1890}, {13'sd2157, 9'sd201, 11'sd-846}, {13'sd3102, 12'sd-1896, 12'sd1575}},
{{10'sd320, 11'sd-537, 12'sd1552}, {14'sd5025, 12'sd-1183, 10'sd-398}, {12'sd1617, 11'sd792, 11'sd-552}},
{{12'sd-1326, 13'sd2403, 13'sd-3441}, {13'sd-2208, 12'sd-1597, 13'sd-3015}, {11'sd641, 12'sd-2016, 12'sd-1346}},
{{13'sd2093, 12'sd1520, 11'sd699}, {12'sd-2018, 12'sd1851, 13'sd2663}, {13'sd-2651, 12'sd-1992, 12'sd1260}},
{{13'sd-2605, 11'sd-584, 12'sd1413}, {14'sd-5333, 12'sd-1806, 10'sd-462}, {14'sd-5442, 14'sd-5554, 12'sd-1412}},
{{13'sd2299, 12'sd1958, 12'sd-1555}, {7'sd54, 13'sd-3516, 11'sd736}, {14'sd4124, 12'sd1843, 12'sd1714}},
{{14'sd-4465, 12'sd-1205, 12'sd-1029}, {13'sd2925, 9'sd187, 13'sd3447}, {12'sd-1386, 8'sd114, 12'sd1675}},
{{13'sd2570, 13'sd-2195, 12'sd1086}, {13'sd3793, 12'sd1767, 10'sd384}, {13'sd3280, 12'sd1188, 10'sd478}},
{{12'sd-1665, 11'sd-614, 13'sd3368}, {13'sd2682, 12'sd-1126, 12'sd1285}, {12'sd1362, 12'sd1888, 13'sd2962}}},
{
{{12'sd-1689, 10'sd-283, 12'sd1564}, {12'sd1806, 12'sd-1177, 12'sd-1514}, {12'sd1246, 11'sd-523, 11'sd-699}},
{{12'sd1796, 13'sd-2450, 10'sd-319}, {13'sd-2620, 13'sd2050, 13'sd-2258}, {11'sd913, 12'sd-1929, 12'sd-1543}},
{{13'sd2375, 10'sd-422, 10'sd-455}, {11'sd585, 11'sd648, 13'sd2471}, {13'sd2499, 11'sd660, 9'sd132}},
{{9'sd-179, 12'sd1486, 13'sd2387}, {12'sd-1228, 12'sd-1260, 12'sd-1277}, {13'sd-2098, 10'sd-343, 4'sd6}},
{{11'sd845, 13'sd2097, 11'sd-603}, {12'sd1794, 11'sd952, 12'sd1247}, {13'sd2942, 14'sd4168, 12'sd1517}},
{{11'sd780, 9'sd165, 14'sd-4196}, {12'sd1714, 10'sd393, 13'sd-2093}, {12'sd-1477, 12'sd1699, 13'sd-3304}},
{{10'sd-302, 13'sd2519, 12'sd1179}, {8'sd-102, 13'sd-2143, 13'sd2073}, {13'sd2953, 11'sd-871, 12'sd1499}},
{{11'sd531, 11'sd-522, 12'sd-1381}, {12'sd1567, 11'sd-815, 11'sd-1013}, {9'sd-196, 11'sd910, 12'sd-1939}},
{{12'sd1740, 12'sd1921, 12'sd2025}, {13'sd2369, 7'sd-50, 9'sd-168}, {11'sd575, 12'sd-1574, 13'sd2475}},
{{11'sd-638, 13'sd3248, 11'sd-974}, {13'sd2351, 10'sd296, 13'sd2394}, {12'sd-1840, 12'sd1895, 13'sd-2157}},
{{12'sd1099, 10'sd395, 13'sd2952}, {12'sd1510, 13'sd3014, 12'sd1487}, {11'sd-623, 10'sd310, 5'sd10}},
{{12'sd-1962, 10'sd452, 13'sd-2735}, {13'sd2336, 12'sd1037, 13'sd-2431}, {12'sd1409, 12'sd-2002, 13'sd-2321}},
{{11'sd759, 11'sd634, 12'sd-1427}, {11'sd629, 13'sd3088, 12'sd-1200}, {12'sd1807, 12'sd1470, 10'sd318}},
{{11'sd-977, 12'sd1223, 13'sd-2364}, {12'sd2024, 10'sd478, 11'sd-856}, {12'sd1832, 10'sd348, 11'sd688}},
{{12'sd1097, 13'sd3540, 13'sd2289}, {9'sd-169, 13'sd3690, 8'sd-86}, {7'sd-49, 10'sd500, 11'sd568}},
{{12'sd2037, 12'sd-1957, 12'sd-1510}, {13'sd2119, 12'sd1870, 12'sd1526}, {11'sd851, 12'sd-1529, 12'sd-1556}},
{{13'sd-2048, 11'sd-719, 11'sd1011}, {13'sd-2859, 9'sd-160, 12'sd-1136}, {11'sd-714, 12'sd2015, 13'sd2118}},
{{13'sd3073, 12'sd-1192, 8'sd118}, {8'sd68, 11'sd-985, 12'sd1569}, {12'sd1478, 11'sd595, 13'sd2529}},
{{12'sd-1536, 11'sd968, 13'sd2305}, {12'sd-1710, 12'sd-1088, 11'sd-993}, {13'sd2364, 12'sd-1180, 12'sd1515}},
{{11'sd839, 11'sd936, 12'sd1870}, {12'sd-1201, 10'sd-333, 13'sd-2750}, {10'sd278, 12'sd1689, 13'sd2165}},
{{8'sd92, 8'sd80, 8'sd-110}, {13'sd-2278, 13'sd2384, 11'sd693}, {13'sd-2175, 13'sd-2470, 11'sd-636}},
{{11'sd762, 13'sd-2869, 13'sd-2739}, {11'sd-728, 12'sd-2004, 12'sd1901}, {12'sd-1885, 12'sd1360, 13'sd-2694}},
{{13'sd-2280, 12'sd1994, 9'sd-179}, {8'sd-67, 13'sd2381, 12'sd1561}, {13'sd2273, 9'sd-251, 7'sd-51}},
{{12'sd-1572, 12'sd-1938, 11'sd-625}, {12'sd1793, 10'sd480, 12'sd1974}, {12'sd-1027, 11'sd881, 13'sd2489}},
{{12'sd1984, 12'sd1835, 12'sd1235}, {12'sd-2035, 11'sd-930, 12'sd-1345}, {11'sd-947, 12'sd-1970, 13'sd-2188}},
{{13'sd2977, 12'sd1915, 11'sd-983}, {13'sd2676, 13'sd-2067, 13'sd2363}, {7'sd63, 13'sd2252, 11'sd532}},
{{13'sd2416, 12'sd1099, 13'sd2313}, {13'sd2579, 11'sd-586, 12'sd1670}, {14'sd4865, 13'sd2523, 8'sd106}},
{{13'sd2633, 11'sd-933, 12'sd-1454}, {13'sd2949, 11'sd-1008, 11'sd-544}, {12'sd-1051, 10'sd503, 10'sd450}},
{{9'sd-189, 12'sd1203, 13'sd-2319}, {12'sd-1296, 5'sd14, 12'sd1263}, {12'sd-1634, 13'sd2140, 10'sd408}},
{{12'sd1439, 13'sd2127, 12'sd-1661}, {13'sd-2127, 13'sd2349, 13'sd-2223}, {10'sd307, 13'sd-2166, 12'sd-1686}},
{{12'sd-1801, 11'sd553, 10'sd-481}, {10'sd-408, 12'sd1033, 11'sd-603}, {12'sd-1283, 13'sd2125, 9'sd187}},
{{12'sd1651, 12'sd-1723, 12'sd1733}, {12'sd-1262, 12'sd1133, 13'sd2127}, {13'sd2482, 9'sd-163, 10'sd-461}},
{{11'sd597, 12'sd-1693, 12'sd2018}, {12'sd1374, 13'sd-2589, 13'sd2153}, {12'sd-2022, 12'sd1584, 13'sd2107}},
{{9'sd251, 11'sd983, 12'sd2041}, {13'sd-2525, 13'sd-2329, 13'sd-2558}, {12'sd-1314, 12'sd1927, 11'sd-755}},
{{13'sd-2667, 10'sd476, 13'sd-2134}, {11'sd-624, 11'sd-713, 12'sd1505}, {11'sd-864, 12'sd-1568, 13'sd-2252}},
{{12'sd-1064, 13'sd-2699, 12'sd-1657}, {10'sd438, 12'sd-1483, 10'sd329}, {11'sd-918, 12'sd1773, 12'sd2011}},
{{12'sd1024, 1'sd0, 12'sd1249}, {12'sd1050, 10'sd366, 7'sd-48}, {9'sd204, 8'sd-65, 11'sd-802}},
{{13'sd2106, 12'sd1777, 13'sd-2156}, {12'sd1954, 11'sd-512, 13'sd2787}, {13'sd2884, 9'sd-167, 13'sd2084}},
{{12'sd1651, 9'sd-128, 10'sd-507}, {11'sd788, 12'sd1573, 12'sd-1561}, {12'sd1134, 12'sd1727, 12'sd-1420}},
{{11'sd-905, 11'sd577, 11'sd981}, {11'sd869, 12'sd1177, 13'sd2763}, {12'sd-1727, 13'sd-2589, 12'sd1065}},
{{11'sd729, 12'sd-1861, 11'sd-886}, {9'sd-170, 10'sd-484, 12'sd-1416}, {6'sd-16, 13'sd2632, 13'sd2413}},
{{12'sd1460, 13'sd-2055, 12'sd1307}, {13'sd2273, 13'sd2078, 13'sd2527}, {11'sd859, 11'sd577, 10'sd449}},
{{13'sd2403, 13'sd2670, 11'sd-615}, {12'sd-1213, 13'sd2058, 13'sd2077}, {9'sd196, 11'sd607, 13'sd2620}},
{{13'sd2212, 10'sd-436, 11'sd-572}, {11'sd793, 13'sd3458, 13'sd-2078}, {12'sd1936, 13'sd3687, 12'sd-2039}},
{{12'sd-1483, 13'sd2280, 11'sd-556}, {12'sd-1258, 13'sd-2376, 12'sd1320}, {11'sd861, 12'sd1343, 13'sd-2656}},
{{11'sd-524, 13'sd-2591, 12'sd-2025}, {13'sd-2736, 13'sd-2285, 12'sd-1198}, {13'sd2117, 13'sd-2291, 12'sd1753}},
{{10'sd-384, 12'sd1077, 7'sd-62}, {12'sd1915, 12'sd1136, 13'sd-3051}, {13'sd2177, 13'sd-2051, 13'sd-2895}},
{{11'sd756, 13'sd2927, 10'sd483}, {13'sd3348, 10'sd-329, 12'sd-1805}, {12'sd1602, 12'sd-1542, 13'sd2935}},
{{10'sd-416, 9'sd169, 13'sd-3346}, {13'sd2470, 13'sd-2964, 13'sd-2810}, {11'sd-775, 13'sd-2996, 11'sd-667}},
{{11'sd571, 12'sd1398, 12'sd-1302}, {13'sd-3191, 13'sd-3473, 12'sd1209}, {8'sd126, 10'sd-487, 13'sd-2625}},
{{11'sd744, 12'sd-1964, 11'sd788}, {12'sd1360, 12'sd1659, 12'sd-1147}, {12'sd1194, 13'sd-2327, 13'sd2394}},
{{11'sd-658, 13'sd-2239, 12'sd-1965}, {11'sd-923, 12'sd-1762, 11'sd-614}, {12'sd-1155, 12'sd1322, 11'sd696}},
{{11'sd-760, 10'sd411, 12'sd-1061}, {13'sd-2285, 10'sd-273, 11'sd-687}, {12'sd1168, 12'sd-1841, 13'sd-2267}},
{{8'sd107, 12'sd-1096, 11'sd853}, {12'sd1183, 10'sd258, 13'sd-2105}, {12'sd1736, 12'sd1938, 12'sd-1289}},
{{12'sd1742, 13'sd2874, 13'sd3658}, {12'sd1232, 12'sd1913, 12'sd1994}, {12'sd-1349, 12'sd-1287, 10'sd360}},
{{12'sd1425, 12'sd-1433, 12'sd-1897}, {13'sd-2357, 11'sd-813, 12'sd-1405}, {11'sd-561, 10'sd299, 12'sd-1785}},
{{13'sd2872, 12'sd1061, 11'sd977}, {11'sd-756, 13'sd3208, 13'sd4080}, {13'sd2281, 9'sd143, 13'sd3954}},
{{12'sd-1372, 11'sd-897, 12'sd-1668}, {13'sd2421, 12'sd1329, 13'sd2684}, {12'sd-1257, 13'sd2267, 13'sd2297}},
{{12'sd1420, 10'sd303, 11'sd929}, {13'sd-2192, 12'sd-1472, 13'sd2481}, {12'sd1975, 12'sd-1944, 11'sd533}},
{{10'sd483, 11'sd589, 11'sd594}, {12'sd-1357, 11'sd-737, 13'sd-2103}, {6'sd-18, 11'sd870, 10'sd-509}},
{{8'sd69, 12'sd-1251, 13'sd-2450}, {8'sd-121, 11'sd-979, 13'sd2168}, {12'sd-1721, 8'sd-99, 13'sd-2243}},
{{12'sd1149, 9'sd-179, 12'sd-1947}, {12'sd-1678, 10'sd273, 12'sd1674}, {11'sd620, 13'sd2583, 9'sd214}},
{{11'sd989, 13'sd-2149, 12'sd1681}, {7'sd49, 13'sd-2119, 8'sd-66}, {12'sd-1351, 12'sd1247, 11'sd-669}},
{{9'sd-203, 11'sd-834, 12'sd-1361}, {12'sd1434, 10'sd301, 12'sd1407}, {12'sd1562, 13'sd2487, 13'sd-2864}}},
{
{{11'sd-532, 13'sd-2373, 10'sd-259}, {10'sd302, 13'sd2509, 12'sd-1286}, {9'sd-158, 12'sd1990, 13'sd2402}},
{{9'sd-205, 12'sd1307, 12'sd1615}, {12'sd-2023, 12'sd1163, 13'sd2391}, {11'sd989, 11'sd675, 12'sd-1318}},
{{13'sd-3198, 12'sd-1581, 13'sd-2359}, {11'sd-707, 12'sd1307, 13'sd-2582}, {11'sd-814, 11'sd-860, 13'sd2738}},
{{12'sd-1525, 11'sd839, 13'sd-2252}, {11'sd-817, 12'sd-1589, 12'sd-1080}, {12'sd-1186, 9'sd132, 10'sd339}},
{{11'sd881, 12'sd-1228, 10'sd-267}, {13'sd2288, 10'sd348, 13'sd2785}, {12'sd1100, 13'sd3890, 13'sd3379}},
{{11'sd-630, 13'sd-2441, 12'sd-1600}, {10'sd282, 13'sd-2831, 11'sd1014}, {13'sd-2670, 9'sd232, 11'sd-630}},
{{11'sd-948, 12'sd1052, 10'sd370}, {13'sd3893, 13'sd-2175, 13'sd2686}, {10'sd412, 12'sd-1274, 10'sd-460}},
{{12'sd-1145, 13'sd2409, 13'sd-2702}, {13'sd2111, 12'sd1642, 12'sd1633}, {12'sd-1902, 12'sd-1578, 8'sd-92}},
{{8'sd88, 8'sd-71, 13'sd-2154}, {11'sd-638, 12'sd1146, 12'sd1438}, {10'sd-447, 13'sd2932, 12'sd-1666}},
{{12'sd-1534, 12'sd1124, 7'sd42}, {9'sd-172, 10'sd-461, 12'sd1366}, {12'sd1806, 13'sd-2739, 12'sd1643}},
{{13'sd-2430, 12'sd1156, 12'sd-1649}, {12'sd-1786, 12'sd-1632, 11'sd731}, {12'sd1625, 13'sd2088, 10'sd477}},
{{7'sd-41, 7'sd-58, 12'sd-1230}, {13'sd-2558, 12'sd1833, 12'sd1605}, {10'sd-274, 13'sd-2406, 12'sd1509}},
{{13'sd2092, 10'sd330, 8'sd-94}, {13'sd2220, 13'sd2426, 12'sd-1339}, {12'sd-1470, 11'sd794, 11'sd756}},
{{12'sd-1393, 12'sd1552, 12'sd1970}, {7'sd-33, 12'sd-1883, 7'sd35}, {12'sd-1922, 12'sd-1248, 13'sd-2899}},
{{12'sd1911, 12'sd1946, 12'sd1221}, {10'sd446, 7'sd63, 12'sd1942}, {11'sd552, 11'sd-805, 13'sd2246}},
{{9'sd175, 12'sd-1325, 11'sd903}, {13'sd2113, 13'sd-2095, 12'sd-1305}, {12'sd-1817, 11'sd-837, 12'sd2034}},
{{12'sd1257, 12'sd-1940, 12'sd-1265}, {13'sd-2502, 12'sd1828, 9'sd179}, {8'sd-71, 13'sd-2484, 12'sd-1378}},
{{12'sd-1540, 11'sd720, 9'sd137}, {13'sd2871, 11'sd-971, 13'sd2709}, {10'sd386, 11'sd-911, 13'sd2196}},
{{8'sd124, 9'sd241, 13'sd2419}, {12'sd-1673, 13'sd-2606, 10'sd-459}, {13'sd2636, 13'sd-2711, 11'sd688}},
{{13'sd2369, 13'sd2322, 9'sd237}, {10'sd-416, 12'sd1562, 13'sd-2517}, {10'sd314, 12'sd1473, 12'sd1804}},
{{12'sd1509, 12'sd-1280, 10'sd388}, {13'sd2378, 12'sd1464, 12'sd-1608}, {10'sd-396, 12'sd1073, 10'sd-302}},
{{13'sd2759, 12'sd-1369, 10'sd316}, {9'sd-203, 12'sd1902, 11'sd905}, {12'sd-1751, 12'sd-1843, 8'sd-120}},
{{12'sd-1468, 12'sd-1177, 10'sd-506}, {11'sd808, 11'sd542, 11'sd559}, {13'sd2718, 13'sd2843, 12'sd1374}},
{{13'sd2513, 12'sd1749, 12'sd1768}, {10'sd-369, 13'sd2389, 10'sd393}, {8'sd93, 13'sd-2667, 6'sd17}},
{{12'sd-1999, 12'sd-1697, 11'sd-546}, {12'sd-1966, 12'sd1494, 10'sd411}, {10'sd-329, 12'sd-2000, 12'sd1814}},
{{7'sd58, 10'sd-299, 13'sd2589}, {13'sd2682, 12'sd1256, 11'sd-710}, {11'sd1023, 13'sd2987, 13'sd2415}},
{{12'sd-1357, 12'sd-1516, 13'sd-3758}, {12'sd-1856, 13'sd-2951, 10'sd338}, {12'sd-1737, 11'sd977, 11'sd-761}},
{{10'sd-260, 10'sd408, 13'sd-2051}, {11'sd-985, 13'sd2348, 13'sd2710}, {11'sd893, 13'sd2130, 12'sd1464}},
{{10'sd-452, 13'sd-2140, 11'sd-639}, {12'sd2034, 12'sd1948, 11'sd865}, {12'sd1261, 12'sd1703, 11'sd-691}},
{{12'sd-1487, 13'sd-2382, 11'sd725}, {7'sd49, 7'sd44, 13'sd-3095}, {12'sd-1691, 12'sd-1760, 12'sd1186}},
{{12'sd-1748, 11'sd-827, 13'sd-2542}, {9'sd157, 12'sd1921, 13'sd2111}, {13'sd-2169, 10'sd-266, 13'sd2542}},
{{12'sd-1805, 12'sd-1219, 12'sd-1798}, {10'sd370, 13'sd2208, 11'sd965}, {12'sd1422, 11'sd799, 12'sd1142}},
{{12'sd-2010, 10'sd381, 12'sd1535}, {10'sd480, 12'sd-1991, 11'sd857}, {12'sd-1533, 13'sd2425, 9'sd151}},
{{12'sd1606, 12'sd1566, 9'sd-183}, {12'sd1502, 9'sd227, 8'sd81}, {10'sd418, 10'sd309, 12'sd-1550}},
{{11'sd-590, 12'sd-1301, 8'sd76}, {12'sd1646, 13'sd-3334, 13'sd-2752}, {11'sd-671, 8'sd-125, 7'sd-32}},
{{12'sd-1359, 13'sd3124, 12'sd1443}, {10'sd479, 13'sd3064, 12'sd1574}, {12'sd1657, 12'sd-1710, 13'sd-2803}},
{{12'sd1313, 13'sd-3491, 12'sd-1106}, {8'sd104, 13'sd-2801, 13'sd-2630}, {12'sd1657, 13'sd-2679, 13'sd-3847}},
{{11'sd-552, 9'sd-165, 12'sd-1570}, {11'sd-927, 12'sd-1760, 12'sd-1297}, {13'sd2900, 13'sd2104, 10'sd-342}},
{{13'sd2435, 12'sd-1575, 12'sd2040}, {11'sd-667, 13'sd-2206, 12'sd1361}, {12'sd-1787, 12'sd-1927, 12'sd1987}},
{{13'sd-2852, 13'sd2415, 13'sd-2531}, {12'sd1548, 11'sd980, 13'sd-2255}, {13'sd-2148, 9'sd180, 13'sd2255}},
{{12'sd2026, 12'sd1138, 12'sd1938}, {11'sd669, 12'sd-1262, 12'sd1368}, {12'sd1901, 12'sd1331, 12'sd1986}},
{{12'sd1411, 13'sd2341, 12'sd1296}, {10'sd458, 11'sd989, 12'sd1973}, {12'sd-1165, 13'sd2451, 11'sd640}},
{{12'sd-1310, 11'sd-718, 12'sd-1834}, {11'sd885, 13'sd-2406, 12'sd-1086}, {13'sd-3326, 12'sd1375, 12'sd-1232}},
{{13'sd-2263, 14'sd-7921, 13'sd-3663}, {12'sd1548, 12'sd-1389, 14'sd-4183}, {12'sd1659, 10'sd-313, 12'sd-1404}},
{{12'sd1334, 12'sd-1248, 10'sd-260}, {10'sd403, 12'sd1177, 12'sd1526}, {12'sd-1078, 12'sd1182, 12'sd1346}},
{{9'sd-168, 12'sd-1984, 12'sd1759}, {13'sd-2678, 11'sd740, 12'sd-1627}, {9'sd-224, 12'sd-1979, 10'sd-300}},
{{10'sd-289, 11'sd-655, 13'sd-2533}, {12'sd-1831, 12'sd-1524, 13'sd-2410}, {10'sd384, 11'sd1012, 12'sd2045}},
{{12'sd-1073, 12'sd-1475, 10'sd356}, {9'sd-240, 13'sd-2699, 11'sd1022}, {11'sd-1010, 13'sd3213, 12'sd1062}},
{{14'sd-4128, 9'sd238, 13'sd-3456}, {13'sd-2869, 13'sd-2272, 11'sd-1003}, {13'sd-3534, 11'sd942, 12'sd1238}},
{{13'sd2199, 13'sd2540, 10'sd499}, {11'sd696, 9'sd150, 11'sd-986}, {12'sd1402, 11'sd615, 13'sd3106}},
{{12'sd1229, 10'sd-387, 9'sd-253}, {12'sd-1053, 11'sd694, 11'sd-560}, {12'sd1632, 9'sd-235, 13'sd2414}},
{{9'sd-199, 11'sd1005, 13'sd2718}, {10'sd395, 12'sd1797, 12'sd-1363}, {9'sd206, 12'sd-1920, 12'sd1127}},
{{11'sd589, 11'sd765, 6'sd17}, {12'sd-2013, 12'sd1563, 8'sd116}, {11'sd1006, 13'sd2810, 11'sd-518}},
{{8'sd-65, 13'sd2576, 12'sd-1030}, {12'sd-1263, 13'sd-2243, 13'sd-2816}, {12'sd1320, 12'sd-2002, 12'sd1774}},
{{12'sd1384, 13'sd2424, 11'sd-834}, {8'sd104, 10'sd-298, 11'sd-817}, {10'sd318, 9'sd213, 13'sd3156}},
{{13'sd-2733, 12'sd-1784, 9'sd136}, {12'sd1901, 11'sd537, 13'sd-2135}, {12'sd1397, 11'sd-783, 12'sd1600}},
{{14'sd5144, 12'sd1107, 13'sd2391}, {14'sd5550, 11'sd913, 13'sd2882}, {7'sd-46, 13'sd2480, 11'sd-949}},
{{13'sd-2668, 12'sd1724, 13'sd-2269}, {12'sd-1811, 9'sd182, 12'sd1918}, {12'sd1331, 13'sd3437, 13'sd2735}},
{{10'sd312, 6'sd-24, 12'sd-1513}, {11'sd-947, 12'sd1374, 12'sd1193}, {12'sd-1653, 11'sd-946, 12'sd-1543}},
{{12'sd-1900, 12'sd-1411, 13'sd3505}, {12'sd-1424, 10'sd373, 13'sd2985}, {13'sd-3036, 13'sd2156, 13'sd2702}},
{{11'sd-581, 12'sd1884, 12'sd-2019}, {13'sd2341, 8'sd-84, 11'sd523}, {11'sd-736, 10'sd416, 12'sd-1442}},
{{13'sd2612, 10'sd-369, 9'sd-148}, {12'sd-2011, 12'sd-1223, 12'sd-1292}, {12'sd-1378, 12'sd1114, 13'sd2965}},
{{12'sd1117, 13'sd-2904, 9'sd-160}, {13'sd-2539, 12'sd-1992, 12'sd1572}, {12'sd-1310, 12'sd1061, 13'sd-2048}},
{{12'sd-1279, 12'sd1164, 10'sd488}, {10'sd-331, 13'sd-2841, 12'sd-1476}, {12'sd1181, 12'sd1191, 13'sd-3227}}},
{
{{12'sd-1382, 10'sd345, 12'sd1867}, {11'sd933, 10'sd-271, 13'sd-2232}, {10'sd444, 11'sd599, 11'sd669}},
{{11'sd948, 13'sd2635, 10'sd460}, {12'sd-1609, 12'sd1472, 12'sd1702}, {13'sd-2080, 12'sd-1907, 13'sd2139}},
{{12'sd-1506, 11'sd942, 11'sd674}, {12'sd1875, 12'sd-1818, 11'sd965}, {10'sd-395, 13'sd2081, 12'sd-1804}},
{{11'sd863, 12'sd-2000, 5'sd-11}, {12'sd-1100, 8'sd-125, 11'sd654}, {12'sd-1351, 12'sd-1690, 12'sd1449}},
{{13'sd3108, 10'sd-478, 13'sd2738}, {13'sd3421, 12'sd-1377, 11'sd-844}, {12'sd-1159, 11'sd628, 10'sd-330}},
{{11'sd677, 12'sd-1713, 10'sd499}, {12'sd-1232, 13'sd-2618, 13'sd-3554}, {13'sd-2376, 13'sd2305, 12'sd1228}},
{{11'sd752, 12'sd1208, 12'sd1369}, {13'sd2875, 13'sd2829, 11'sd645}, {13'sd2527, 12'sd-1092, 12'sd1841}},
{{12'sd1802, 13'sd-2573, 11'sd790}, {10'sd-451, 13'sd2780, 12'sd-1606}, {11'sd-562, 12'sd-1941, 11'sd787}},
{{12'sd-1543, 13'sd2809, 10'sd509}, {12'sd-1704, 9'sd-227, 12'sd-1595}, {7'sd-49, 12'sd-1540, 11'sd-896}},
{{12'sd-1123, 12'sd-1170, 12'sd-1431}, {11'sd-544, 12'sd-1242, 10'sd483}, {13'sd2392, 9'sd-130, 11'sd572}},
{{12'sd-1094, 11'sd-838, 10'sd-324}, {12'sd-1837, 9'sd-182, 13'sd-2287}, {7'sd-49, 13'sd2289, 13'sd-2789}},
{{9'sd243, 12'sd1555, 8'sd120}, {11'sd728, 12'sd-1978, 12'sd-1047}, {12'sd-1892, 11'sd-813, 12'sd-1727}},
{{12'sd2007, 13'sd2739, 11'sd-561}, {12'sd-1781, 12'sd2016, 12'sd-1780}, {12'sd-1834, 11'sd-912, 12'sd-1370}},
{{9'sd-248, 11'sd-837, 12'sd-1889}, {11'sd780, 10'sd-456, 10'sd383}, {12'sd-1801, 11'sd-982, 12'sd1990}},
{{11'sd659, 12'sd-1820, 12'sd-1154}, {13'sd2053, 12'sd-1618, 13'sd2629}, {11'sd-554, 12'sd1946, 12'sd-1373}},
{{13'sd2772, 12'sd-1638, 12'sd1932}, {13'sd2172, 12'sd1660, 10'sd-265}, {11'sd621, 13'sd-2296, 7'sd-51}},
{{13'sd2272, 13'sd-2069, 13'sd-2575}, {10'sd-452, 12'sd1982, 10'sd-257}, {12'sd-1778, 10'sd-266, 9'sd133}},
{{13'sd3412, 10'sd-489, 12'sd-1151}, {12'sd1813, 13'sd2391, 12'sd-1579}, {11'sd-1002, 13'sd2606, 12'sd1551}},
{{13'sd2625, 13'sd-2453, 13'sd2201}, {12'sd-1458, 9'sd184, 12'sd1857}, {13'sd-2157, 10'sd324, 12'sd1433}},
{{13'sd-2680, 12'sd1665, 13'sd-2400}, {10'sd486, 13'sd2575, 12'sd-1398}, {12'sd-1760, 13'sd-2520, 10'sd-376}},
{{11'sd-902, 12'sd-1458, 10'sd-509}, {10'sd349, 13'sd2241, 12'sd1237}, {2'sd1, 12'sd-1533, 12'sd-1221}},
{{12'sd-1673, 13'sd-2439, 10'sd-294}, {13'sd2613, 12'sd-1039, 11'sd-968}, {12'sd-1050, 12'sd-1273, 13'sd2254}},
{{11'sd898, 12'sd1409, 10'sd-297}, {13'sd-2554, 12'sd1367, 12'sd1734}, {12'sd-2022, 10'sd369, 11'sd-974}},
{{13'sd2525, 13'sd-2782, 12'sd-1216}, {13'sd-2458, 13'sd-2524, 11'sd838}, {11'sd966, 10'sd-470, 13'sd2483}},
{{13'sd2516, 12'sd-1667, 11'sd-895}, {12'sd1819, 12'sd1255, 10'sd338}, {11'sd752, 13'sd2147, 12'sd-1982}},
{{12'sd1346, 10'sd-261, 11'sd581}, {13'sd-2219, 13'sd2642, 11'sd-936}, {10'sd-386, 12'sd1095, 10'sd494}},
{{11'sd987, 13'sd2416, 12'sd-1436}, {13'sd3545, 13'sd3221, 11'sd1017}, {12'sd1303, 11'sd728, 11'sd733}},
{{13'sd2484, 11'sd889, 9'sd-175}, {11'sd581, 5'sd8, 13'sd2244}, {11'sd576, 12'sd1538, 12'sd-1140}},
{{12'sd1286, 12'sd1235, 10'sd264}, {10'sd-316, 12'sd-1701, 11'sd-723}, {12'sd1245, 10'sd-452, 9'sd196}},
{{9'sd-149, 10'sd-356, 13'sd-2094}, {9'sd-183, 13'sd2334, 13'sd-2741}, {12'sd1967, 13'sd-2895, 13'sd2597}},
{{11'sd-740, 13'sd-2860, 12'sd1718}, {13'sd2301, 13'sd2435, 7'sd45}, {8'sd76, 12'sd1640, 11'sd-865}},
{{11'sd-675, 12'sd1051, 12'sd1048}, {11'sd-536, 12'sd-1704, 12'sd-1579}, {13'sd2342, 13'sd-2084, 11'sd878}},
{{13'sd-2223, 8'sd-100, 12'sd1143}, {13'sd-2324, 10'sd335, 12'sd1477}, {13'sd2298, 13'sd-2285, 11'sd-726}},
{{13'sd3425, 12'sd1674, 13'sd-2351}, {11'sd-905, 12'sd1426, 13'sd2345}, {10'sd402, 13'sd2558, 10'sd469}},
{{10'sd272, 12'sd1971, 13'sd3017}, {12'sd-1776, 13'sd-2138, 12'sd-1504}, {10'sd-326, 12'sd-1573, 13'sd2330}},
{{12'sd1823, 13'sd-2385, 10'sd-299}, {11'sd-898, 7'sd56, 11'sd-907}, {12'sd1375, 13'sd2798, 12'sd1250}},
{{11'sd680, 14'sd-4901, 13'sd-2942}, {13'sd2217, 12'sd-1728, 12'sd1147}, {10'sd-274, 13'sd-2904, 13'sd-2644}},
{{11'sd-736, 4'sd-6, 11'sd-619}, {10'sd492, 12'sd1311, 12'sd2040}, {10'sd505, 12'sd1208, 13'sd3101}},
{{10'sd476, 12'sd-1855, 13'sd2974}, {11'sd1022, 13'sd2108, 13'sd-2331}, {12'sd1380, 11'sd863, 13'sd2854}},
{{13'sd2376, 7'sd33, 11'sd-716}, {13'sd2129, 12'sd1040, 12'sd1477}, {12'sd1778, 11'sd-907, 12'sd-1569}},
{{13'sd2582, 12'sd1848, 13'sd2781}, {12'sd1073, 13'sd2332, 10'sd-433}, {10'sd384, 9'sd-206, 13'sd2061}},
{{10'sd-322, 9'sd-150, 13'sd-2446}, {11'sd-676, 12'sd1752, 12'sd1292}, {10'sd492, 13'sd-2581, 12'sd1554}},
{{12'sd-1099, 11'sd539, 13'sd2546}, {13'sd3202, 13'sd3057, 11'sd792}, {13'sd2565, 12'sd1221, 12'sd1101}},
{{13'sd-2636, 12'sd1210, 11'sd-604}, {12'sd1547, 13'sd2658, 13'sd2304}, {13'sd2733, 13'sd2229, 11'sd819}},
{{12'sd-1245, 10'sd433, 11'sd-817}, {9'sd171, 9'sd-128, 12'sd2021}, {12'sd1182, 12'sd-1255, 12'sd-1380}},
{{11'sd-945, 13'sd-3052, 13'sd-2218}, {12'sd1288, 12'sd1344, 13'sd-2507}, {11'sd-541, 9'sd-173, 6'sd-29}},
{{10'sd-401, 13'sd2507, 9'sd-138}, {7'sd-40, 10'sd479, 10'sd288}, {8'sd-64, 13'sd2204, 13'sd-2130}},
{{12'sd-1441, 12'sd-1218, 11'sd761}, {10'sd-508, 13'sd-2231, 11'sd-523}, {13'sd3384, 13'sd-2124, 10'sd-503}},
{{8'sd66, 13'sd-2484, 12'sd-1989}, {12'sd1851, 13'sd-2595, 12'sd-1278}, {13'sd2512, 11'sd862, 12'sd1257}},
{{12'sd-1649, 9'sd221, 12'sd1678}, {12'sd1792, 13'sd-2337, 12'sd-1745}, {12'sd1401, 12'sd-1940, 13'sd-2833}},
{{13'sd2543, 12'sd1843, 12'sd-1125}, {13'sd2639, 10'sd468, 13'sd2441}, {13'sd-2106, 13'sd2205, 13'sd3057}},
{{13'sd-2365, 13'sd-2171, 12'sd-1984}, {13'sd2338, 13'sd-2858, 12'sd1951}, {12'sd1586, 10'sd-461, 11'sd544}},
{{12'sd-1198, 11'sd966, 12'sd-1099}, {11'sd-686, 11'sd852, 11'sd-865}, {13'sd-2761, 11'sd708, 11'sd824}},
{{13'sd-2060, 8'sd-82, 12'sd1458}, {12'sd-2010, 11'sd718, 12'sd-1993}, {12'sd-1795, 11'sd-588, 10'sd-363}},
{{12'sd1424, 11'sd521, 10'sd511}, {6'sd-20, 10'sd-445, 12'sd-1766}, {11'sd939, 13'sd2901, 13'sd2346}},
{{13'sd-3028, 11'sd991, 13'sd-2549}, {12'sd1559, 12'sd-1289, 6'sd20}, {13'sd2480, 13'sd-2531, 11'sd-570}},
{{12'sd-1618, 12'sd1548, 12'sd1683}, {7'sd-41, 12'sd1292, 13'sd2906}, {12'sd-2008, 11'sd-515, 13'sd3406}},
{{12'sd1664, 7'sd-50, 11'sd-740}, {12'sd1884, 11'sd963, 13'sd3040}, {13'sd-2571, 13'sd2151, 13'sd2560}},
{{12'sd2038, 12'sd-1374, 11'sd-725}, {11'sd-617, 12'sd-1772, 12'sd-2027}, {12'sd1296, 13'sd-2799, 11'sd920}},
{{11'sd653, 11'sd654, 12'sd-1098}, {12'sd-1191, 12'sd1308, 13'sd2103}, {13'sd3628, 11'sd930, 11'sd1003}},
{{12'sd-1655, 11'sd839, 12'sd1622}, {11'sd738, 12'sd1389, 12'sd1026}, {9'sd175, 12'sd-1700, 13'sd2998}},
{{8'sd-71, 12'sd1761, 12'sd-1569}, {9'sd161, 12'sd-1162, 9'sd234}, {13'sd-2183, 12'sd-1854, 12'sd1099}},
{{12'sd-1034, 9'sd254, 12'sd-1464}, {12'sd-1286, 8'sd-126, 11'sd746}, {11'sd518, 11'sd-869, 7'sd61}},
{{10'sd-480, 11'sd934, 11'sd-868}, {12'sd-1208, 13'sd2810, 10'sd322}, {12'sd-1516, 12'sd1888, 12'sd-1323}}},
{
{{13'sd2634, 13'sd2853, 11'sd-810}, {13'sd2479, 11'sd-810, 11'sd674}, {10'sd-420, 8'sd71, 13'sd2542}},
{{11'sd732, 13'sd-2534, 13'sd-2226}, {11'sd-654, 12'sd-1618, 13'sd-2099}, {13'sd-2375, 10'sd426, 13'sd2157}},
{{13'sd-2331, 12'sd1847, 12'sd-1627}, {11'sd718, 13'sd-2442, 13'sd2609}, {12'sd-1029, 10'sd-433, 11'sd521}},
{{12'sd1378, 11'sd963, 11'sd588}, {11'sd-628, 12'sd-2013, 13'sd-2120}, {13'sd2387, 11'sd547, 9'sd-148}},
{{14'sd-5458, 12'sd-1448, 11'sd988}, {9'sd-230, 12'sd-1627, 13'sd2155}, {6'sd-17, 12'sd1996, 13'sd3040}},
{{11'sd-894, 9'sd-129, 9'sd-159}, {12'sd1893, 13'sd-2935, 12'sd-1448}, {9'sd210, 10'sd-271, 13'sd-3619}},
{{12'sd1098, 12'sd-1903, 13'sd-2649}, {13'sd-3826, 12'sd-1541, 12'sd-1251}, {10'sd317, 11'sd-855, 8'sd78}},
{{13'sd2979, 11'sd-619, 8'sd-64}, {11'sd836, 12'sd-1386, 12'sd1378}, {11'sd-601, 11'sd1015, 11'sd-774}},
{{11'sd558, 13'sd-2525, 12'sd-1087}, {10'sd-314, 12'sd-1123, 13'sd2819}, {10'sd-488, 13'sd2504, 11'sd-552}},
{{13'sd2340, 13'sd-2793, 3'sd2}, {13'sd2907, 13'sd-2274, 9'sd172}, {12'sd1971, 12'sd-1833, 13'sd2596}},
{{10'sd-482, 12'sd-1306, 10'sd-406}, {11'sd554, 11'sd764, 13'sd-2101}, {12'sd1485, 12'sd1751, 13'sd2116}},
{{12'sd-1727, 13'sd2284, 9'sd139}, {10'sd-262, 13'sd2112, 13'sd3211}, {12'sd-1455, 9'sd168, 11'sd-641}},
{{12'sd1908, 12'sd-1904, 12'sd1923}, {12'sd1565, 10'sd-261, 12'sd1111}, {9'sd-212, 13'sd2492, 12'sd1292}},
{{8'sd89, 13'sd-2363, 11'sd739}, {12'sd-1654, 12'sd-1100, 12'sd-1072}, {13'sd-2761, 13'sd2549, 13'sd-2566}},
{{13'sd-3369, 12'sd-1625, 11'sd942}, {11'sd-569, 12'sd-1322, 12'sd1916}, {13'sd3198, 11'sd876, 12'sd1131}},
{{12'sd1214, 13'sd2641, 9'sd183}, {13'sd2683, 12'sd-1028, 12'sd-1145}, {12'sd-1387, 11'sd-548, 13'sd3448}},
{{12'sd-1815, 13'sd-2186, 12'sd-1553}, {11'sd-724, 11'sd953, 13'sd-2569}, {13'sd-2645, 13'sd-2578, 13'sd-2491}},
{{10'sd-380, 11'sd818, 12'sd1569}, {12'sd-1160, 12'sd-1151, 12'sd-1850}, {13'sd2690, 13'sd2202, 13'sd2287}},
{{12'sd-1566, 13'sd2139, 12'sd1348}, {11'sd592, 11'sd-884, 12'sd-1834}, {13'sd2767, 12'sd1530, 8'sd121}},
{{13'sd2056, 13'sd2170, 4'sd-6}, {11'sd925, 12'sd-1617, 10'sd433}, {12'sd-1553, 12'sd-1975, 11'sd904}},
{{12'sd-1492, 12'sd-1519, 11'sd631}, {9'sd182, 12'sd-1696, 10'sd413}, {11'sd540, 12'sd-1599, 12'sd-1721}},
{{13'sd-2225, 12'sd1356, 11'sd913}, {12'sd2038, 11'sd-874, 13'sd-2791}, {8'sd71, 11'sd-953, 12'sd-1562}},
{{12'sd2004, 11'sd844, 9'sd-153}, {12'sd-1427, 12'sd-1840, 10'sd-276}, {12'sd1154, 13'sd2556, 13'sd2987}},
{{13'sd2097, 11'sd1007, 12'sd1721}, {13'sd2548, 11'sd-626, 13'sd2073}, {8'sd117, 8'sd-99, 13'sd2635}},
{{13'sd2484, 12'sd-1439, 10'sd-326}, {11'sd-722, 11'sd529, 12'sd-1391}, {12'sd2032, 11'sd951, 11'sd-809}},
{{12'sd1032, 12'sd-1413, 12'sd-1937}, {13'sd2604, 13'sd-2676, 12'sd-1469}, {12'sd1271, 8'sd69, 12'sd1993}},
{{7'sd56, 13'sd2224, 10'sd-288}, {12'sd-1088, 13'sd-2178, 12'sd-1344}, {13'sd2455, 12'sd1367, 12'sd1599}},
{{11'sd890, 13'sd-2052, 9'sd164}, {13'sd-2363, 8'sd-78, 11'sd565}, {11'sd-897, 12'sd1934, 13'sd2827}},
{{12'sd-1784, 5'sd8, 7'sd-39}, {11'sd1004, 12'sd1103, 11'sd-797}, {11'sd-684, 12'sd1831, 10'sd-426}},
{{12'sd-1533, 10'sd-282, 12'sd-1258}, {10'sd327, 11'sd-854, 12'sd-1025}, {11'sd953, 13'sd2564, 12'sd-1778}},
{{11'sd-737, 13'sd2204, 11'sd983}, {13'sd2728, 13'sd-2275, 12'sd1279}, {12'sd1604, 12'sd1682, 13'sd-2158}},
{{12'sd-1223, 12'sd-1091, 13'sd2608}, {13'sd-2186, 11'sd-939, 11'sd-856}, {12'sd-1694, 10'sd325, 10'sd352}},
{{11'sd635, 13'sd2723, 10'sd-312}, {10'sd-268, 12'sd1587, 12'sd-1884}, {10'sd421, 12'sd1289, 12'sd1616}},
{{13'sd-2227, 12'sd1479, 11'sd595}, {13'sd-2504, 13'sd2156, 12'sd2021}, {10'sd415, 12'sd1251, 11'sd-797}},
{{12'sd-1860, 11'sd513, 10'sd-427}, {11'sd-615, 12'sd1838, 11'sd-664}, {11'sd-635, 12'sd-1257, 12'sd-1292}},
{{11'sd-897, 10'sd440, 10'sd-324}, {12'sd-1920, 13'sd2392, 11'sd-516}, {10'sd-489, 12'sd-1745, 12'sd1661}},
{{13'sd2547, 14'sd4582, 13'sd3191}, {12'sd1624, 13'sd2212, 12'sd1221}, {6'sd31, 13'sd-2313, 13'sd-2496}},
{{12'sd1182, 9'sd211, 10'sd443}, {10'sd401, 12'sd1596, 13'sd-2979}, {8'sd-98, 10'sd-511, 9'sd-156}},
{{12'sd-1056, 8'sd-106, 10'sd361}, {11'sd-757, 10'sd315, 13'sd-2661}, {13'sd2640, 11'sd-609, 13'sd2642}},
{{11'sd671, 13'sd2075, 10'sd-426}, {11'sd939, 10'sd313, 13'sd2740}, {13'sd-2139, 13'sd2292, 13'sd2072}},
{{12'sd1593, 13'sd-2963, 12'sd1649}, {12'sd1457, 9'sd-220, 13'sd-3000}, {11'sd807, 13'sd-2068, 7'sd52}},
{{12'sd-1292, 12'sd-1798, 12'sd-1593}, {11'sd700, 12'sd1177, 12'sd1421}, {13'sd2647, 13'sd3405, 11'sd976}},
{{12'sd1690, 13'sd-3042, 12'sd-1607}, {10'sd316, 12'sd1554, 13'sd-2302}, {13'sd2118, 13'sd2096, 11'sd-601}},
{{13'sd-2793, 13'sd-3103, 12'sd1645}, {12'sd1846, 11'sd-907, 11'sd-515}, {13'sd-2439, 13'sd2544, 12'sd-1776}},
{{10'sd334, 10'sd286, 9'sd249}, {12'sd1750, 13'sd2139, 11'sd-935}, {10'sd320, 12'sd-1669, 13'sd2576}},
{{13'sd2823, 12'sd-1349, 13'sd2870}, {13'sd-2069, 12'sd1443, 12'sd-1831}, {12'sd1701, 11'sd-752, 10'sd-295}},
{{13'sd-2469, 12'sd-1363, 13'sd3390}, {13'sd-2820, 12'sd1196, 13'sd3416}, {12'sd-1536, 10'sd-351, 13'sd2097}},
{{13'sd-3519, 13'sd-2619, 12'sd1206}, {13'sd-2334, 12'sd1416, 11'sd774}, {12'sd1613, 10'sd305, 13'sd-2055}},
{{10'sd-460, 9'sd128, 8'sd105}, {10'sd350, 13'sd-2844, 11'sd789}, {11'sd593, 11'sd-933, 12'sd-1311}},
{{13'sd2175, 13'sd3263, 13'sd2792}, {8'sd78, 14'sd4474, 11'sd766}, {12'sd1527, 6'sd-30, 12'sd1411}},
{{13'sd-2092, 10'sd504, 13'sd-3303}, {12'sd1992, 12'sd1622, 11'sd-997}, {12'sd-1594, 11'sd1014, 10'sd311}},
{{11'sd-990, 13'sd-2309, 12'sd-1262}, {13'sd-2109, 8'sd-82, 12'sd-1434}, {13'sd-2334, 9'sd-135, 12'sd-2000}},
{{12'sd-1414, 11'sd-668, 10'sd-333}, {13'sd2403, 10'sd-347, 13'sd2441}, {11'sd530, 9'sd-182, 12'sd1039}},
{{11'sd-867, 13'sd2592, 12'sd-2006}, {13'sd3054, 13'sd-2384, 13'sd-2530}, {12'sd1477, 12'sd-1234, 13'sd-2496}},
{{13'sd-2079, 13'sd-2260, 12'sd1224}, {11'sd-867, 12'sd-2044, 10'sd320}, {13'sd2823, 12'sd1596, 12'sd1826}},
{{13'sd3500, 13'sd2585, 11'sd671}, {11'sd734, 11'sd-788, 12'sd1813}, {12'sd-1370, 12'sd-1687, 13'sd-2974}},
{{13'sd-2227, 10'sd-295, 10'sd-281}, {10'sd261, 9'sd-203, 9'sd215}, {11'sd902, 13'sd2625, 13'sd2672}},
{{13'sd-3670, 13'sd-2089, 13'sd-2229}, {12'sd-1611, 12'sd1112, 10'sd352}, {12'sd1705, 13'sd-2265, 12'sd-1502}},
{{12'sd-1675, 12'sd-1676, 13'sd2747}, {12'sd-1399, 10'sd-327, 12'sd1724}, {11'sd654, 13'sd-2193, 12'sd-1499}},
{{11'sd625, 13'sd-2055, 11'sd-973}, {13'sd2498, 8'sd-121, 12'sd-1917}, {14'sd4616, 11'sd623, 13'sd3022}},
{{10'sd318, 12'sd1378, 13'sd-2573}, {11'sd-770, 10'sd353, 10'sd-369}, {12'sd-1563, 13'sd2725, 13'sd2481}},
{{12'sd-1420, 10'sd403, 8'sd72}, {13'sd2277, 12'sd-1857, 12'sd1867}, {12'sd2038, 11'sd657, 12'sd1987}},
{{10'sd412, 12'sd-1223, 13'sd-2652}, {10'sd347, 4'sd6, 9'sd226}, {11'sd-671, 12'sd1040, 11'sd547}},
{{11'sd822, 10'sd-388, 12'sd-1207}, {8'sd-78, 10'sd293, 13'sd-2096}, {12'sd1805, 13'sd-2926, 12'sd1160}}},
{
{{13'sd-2671, 11'sd708, 9'sd-203}, {13'sd2328, 9'sd-243, 11'sd557}, {13'sd2074, 13'sd2730, 12'sd-1670}},
{{12'sd-1285, 13'sd-2187, 11'sd619}, {12'sd-1586, 12'sd1659, 12'sd-1653}, {11'sd902, 12'sd-1064, 9'sd171}},
{{12'sd1863, 11'sd-542, 13'sd-2143}, {12'sd1344, 10'sd-374, 13'sd-2114}, {11'sd-762, 12'sd1564, 10'sd325}},
{{11'sd981, 10'sd283, 12'sd1614}, {13'sd-2919, 12'sd1159, 13'sd-2322}, {13'sd-2831, 11'sd-699, 11'sd-1018}},
{{12'sd-1344, 12'sd-1995, 13'sd2663}, {11'sd-993, 12'sd-1856, 10'sd421}, {11'sd-577, 11'sd-1014, 6'sd-16}},
{{12'sd1938, 11'sd-742, 13'sd2126}, {12'sd1057, 10'sd418, 9'sd-134}, {12'sd1856, 12'sd-1229, 8'sd74}},
{{5'sd15, 13'sd2514, 11'sd863}, {12'sd-1127, 10'sd407, 10'sd286}, {12'sd-1079, 11'sd748, 12'sd1712}},
{{11'sd-512, 13'sd-2266, 13'sd2825}, {12'sd-1059, 9'sd155, 12'sd1998}, {11'sd-873, 12'sd1210, 13'sd2603}},
{{13'sd-2456, 12'sd1378, 12'sd-2020}, {11'sd-674, 12'sd-1379, 10'sd-419}, {11'sd719, 12'sd1295, 10'sd-359}},
{{13'sd-2742, 9'sd-222, 12'sd1543}, {12'sd1028, 13'sd-2553, 11'sd-785}, {10'sd364, 12'sd-1580, 11'sd-978}},
{{13'sd-2834, 11'sd-921, 13'sd2142}, {9'sd-141, 12'sd-1905, 13'sd2330}, {12'sd1681, 11'sd-516, 12'sd-1560}},
{{13'sd-2718, 12'sd-2014, 12'sd-1765}, {11'sd-651, 12'sd1235, 12'sd1979}, {12'sd1544, 13'sd-2230, 12'sd1628}},
{{12'sd-1276, 13'sd2515, 12'sd-1123}, {13'sd3085, 12'sd-1224, 12'sd1686}, {10'sd-345, 12'sd1325, 13'sd2882}},
{{12'sd-1286, 8'sd-81, 9'sd-223}, {12'sd-1948, 10'sd259, 10'sd385}, {12'sd1781, 13'sd2465, 12'sd1136}},
{{12'sd1358, 9'sd-147, 12'sd-1624}, {11'sd-833, 10'sd256, 12'sd-1903}, {13'sd-3535, 13'sd-3733, 13'sd-2660}},
{{11'sd607, 10'sd-370, 8'sd-111}, {12'sd-1431, 13'sd3221, 12'sd-1822}, {11'sd911, 12'sd-1251, 13'sd2277}},
{{13'sd-2326, 11'sd878, 12'sd-1925}, {12'sd1249, 11'sd-823, 13'sd-2405}, {13'sd2209, 12'sd-1079, 10'sd-333}},
{{13'sd3006, 12'sd-1122, 12'sd1923}, {11'sd620, 12'sd1604, 12'sd-1445}, {13'sd2699, 9'sd-237, 11'sd-514}},
{{12'sd-1829, 12'sd-1295, 10'sd417}, {12'sd-1843, 10'sd437, 11'sd-660}, {13'sd-2438, 13'sd-2659, 10'sd-415}},
{{13'sd-2199, 12'sd-1059, 11'sd-1002}, {12'sd1286, 12'sd1925, 10'sd-427}, {13'sd-2198, 12'sd1588, 12'sd1543}},
{{12'sd-1926, 12'sd1441, 12'sd-1255}, {12'sd1865, 11'sd-685, 13'sd-2196}, {12'sd-1456, 13'sd-2837, 9'sd230}},
{{12'sd1213, 12'sd1546, 12'sd-1104}, {11'sd-828, 12'sd-2005, 9'sd210}, {8'sd-81, 12'sd1388, 13'sd2157}},
{{12'sd2047, 12'sd1921, 13'sd3178}, {12'sd1060, 13'sd2458, 11'sd-520}, {12'sd1489, 13'sd2655, 13'sd2195}},
{{13'sd2321, 13'sd2348, 10'sd-269}, {13'sd-2487, 13'sd-2723, 12'sd-1058}, {12'sd1584, 12'sd1449, 12'sd1730}},
{{12'sd1402, 12'sd1942, 12'sd1955}, {13'sd-2157, 12'sd-1170, 12'sd1389}, {11'sd954, 10'sd-263, 11'sd955}},
{{10'sd469, 9'sd-186, 12'sd-1062}, {13'sd2506, 11'sd-1010, 9'sd-193}, {13'sd2729, 12'sd1059, 11'sd553}},
{{13'sd3223, 13'sd2905, 12'sd1782}, {7'sd62, 10'sd-297, 10'sd-280}, {12'sd-1463, 11'sd-574, 12'sd-1575}},
{{12'sd-1190, 10'sd347, 12'sd-2004}, {9'sd144, 12'sd-1506, 12'sd-1738}, {11'sd909, 11'sd-990, 12'sd1825}},
{{11'sd762, 13'sd2118, 13'sd-2155}, {12'sd1527, 13'sd2101, 12'sd-1671}, {11'sd-788, 11'sd-689, 13'sd-2551}},
{{9'sd148, 13'sd-2156, 13'sd-3011}, {13'sd2072, 11'sd942, 12'sd-1042}, {12'sd-1759, 12'sd-1521, 12'sd2041}},
{{12'sd-1899, 12'sd-1688, 11'sd806}, {12'sd1057, 12'sd-1664, 12'sd1417}, {12'sd-2012, 12'sd1655, 11'sd-921}},
{{11'sd859, 12'sd1436, 12'sd-1983}, {12'sd-1394, 13'sd2341, 13'sd2364}, {13'sd-2267, 13'sd-2203, 13'sd-2248}},
{{12'sd1305, 11'sd-956, 13'sd2387}, {11'sd534, 10'sd363, 11'sd759}, {13'sd2102, 12'sd-1324, 12'sd1669}},
{{10'sd410, 11'sd967, 11'sd859}, {12'sd-1332, 11'sd637, 13'sd-2096}, {12'sd1797, 12'sd-1880, 12'sd-1726}},
{{11'sd969, 12'sd-1678, 13'sd-2262}, {11'sd-690, 10'sd-279, 13'sd2647}, {12'sd-1785, 13'sd-2601, 12'sd1607}},
{{12'sd1896, 7'sd-62, 8'sd78}, {13'sd2256, 13'sd2220, 12'sd1592}, {12'sd-1455, 13'sd-2587, 12'sd-1363}},
{{12'sd-1284, 10'sd384, 13'sd2425}, {11'sd696, 11'sd-563, 10'sd-294}, {9'sd-171, 12'sd-1767, 12'sd-1692}},
{{12'sd1526, 12'sd-1247, 12'sd1549}, {13'sd-2381, 9'sd172, 11'sd-855}, {10'sd318, 13'sd2132, 8'sd117}},
{{13'sd-2515, 12'sd1975, 12'sd-1989}, {11'sd924, 13'sd2222, 12'sd1512}, {12'sd1873, 12'sd-1956, 11'sd783}},
{{13'sd-2277, 11'sd-870, 11'sd-606}, {12'sd-1831, 10'sd-264, 11'sd605}, {10'sd-405, 12'sd2008, 10'sd486}},
{{13'sd-3211, 11'sd-627, 12'sd2019}, {12'sd1061, 13'sd2298, 10'sd-414}, {13'sd-2644, 11'sd514, 12'sd-1780}},
{{9'sd203, 13'sd2660, 12'sd1058}, {12'sd1223, 13'sd2452, 13'sd2063}, {12'sd1383, 10'sd390, 13'sd2411}},
{{12'sd-1247, 10'sd383, 12'sd-1324}, {12'sd-2037, 10'sd-459, 11'sd783}, {12'sd1675, 11'sd1018, 12'sd1456}},
{{13'sd2880, 13'sd3167, 11'sd556}, {13'sd3129, 11'sd895, 12'sd1683}, {13'sd3116, 14'sd5804, 14'sd4700}},
{{10'sd266, 7'sd44, 10'sd399}, {11'sd888, 12'sd1991, 13'sd2671}, {12'sd1422, 10'sd-321, 11'sd-651}},
{{11'sd-517, 11'sd911, 11'sd-574}, {13'sd2464, 11'sd639, 13'sd2337}, {8'sd101, 10'sd369, 12'sd-1406}},
{{13'sd2234, 9'sd204, 11'sd778}, {13'sd2703, 11'sd-536, 9'sd129}, {13'sd-2654, 12'sd-1088, 11'sd819}},
{{12'sd-1901, 12'sd1326, 12'sd-1602}, {13'sd2213, 12'sd1373, 12'sd-1126}, {12'sd-1367, 13'sd-2247, 11'sd656}},
{{13'sd-2482, 11'sd-652, 13'sd-2252}, {10'sd507, 10'sd284, 12'sd1447}, {13'sd2058, 9'sd-181, 12'sd-1076}},
{{12'sd1523, 13'sd-2279, 12'sd-1628}, {12'sd1447, 11'sd-976, 13'sd-2839}, {13'sd3058, 12'sd-1273, 13'sd-3750}},
{{13'sd-3020, 12'sd-1105, 10'sd-434}, {13'sd-2396, 13'sd-2501, 12'sd1240}, {13'sd-2425, 13'sd-2193, 12'sd1424}},
{{12'sd-1611, 11'sd604, 12'sd-1502}, {12'sd1334, 10'sd489, 11'sd845}, {13'sd2767, 13'sd2489, 12'sd-2016}},
{{10'sd-452, 12'sd1114, 13'sd2615}, {13'sd2293, 10'sd305, 12'sd1523}, {11'sd-748, 4'sd-4, 13'sd2615}},
{{13'sd2635, 12'sd-1804, 12'sd1247}, {12'sd-1037, 13'sd-2198, 12'sd-1286}, {12'sd-1114, 12'sd1172, 12'sd2038}},
{{11'sd804, 11'sd-798, 12'sd1098}, {12'sd1684, 11'sd694, 12'sd-1329}, {13'sd2346, 12'sd2040, 12'sd-1933}},
{{12'sd-1666, 13'sd2214, 10'sd-317}, {12'sd-1778, 12'sd-1752, 11'sd882}, {13'sd2137, 11'sd-572, 11'sd746}},
{{12'sd-1127, 11'sd-599, 8'sd-99}, {12'sd1354, 11'sd708, 12'sd1752}, {12'sd1563, 11'sd-529, 14'sd4615}},
{{12'sd-1422, 10'sd360, 11'sd893}, {12'sd1664, 13'sd2187, 12'sd1696}, {11'sd903, 11'sd-605, 12'sd1842}},
{{12'sd1465, 11'sd-899, 13'sd-2667}, {10'sd405, 8'sd114, 13'sd2186}, {9'sd222, 12'sd-1289, 13'sd2285}},
{{13'sd-2886, 12'sd-1805, 12'sd-1851}, {13'sd2620, 12'sd-1085, 12'sd-1593}, {10'sd372, 12'sd1129, 13'sd-2847}},
{{10'sd-370, 13'sd-2168, 10'sd-257}, {12'sd1762, 13'sd-2309, 13'sd2596}, {11'sd582, 12'sd1062, 13'sd2616}},
{{11'sd529, 10'sd287, 13'sd-2360}, {11'sd-921, 12'sd1248, 11'sd-799}, {11'sd691, 11'sd595, 13'sd2610}},
{{12'sd-1315, 11'sd907, 7'sd-43}, {13'sd-2755, 11'sd-537, 13'sd2320}, {5'sd-14, 12'sd1711, 12'sd1674}},
{{12'sd2035, 11'sd-524, 11'sd-797}, {12'sd-1981, 12'sd-1774, 13'sd-3186}, {11'sd-941, 12'sd-1475, 13'sd-3232}}}},
// Weights for conv3_weight
{
{
{{11'sd-978, 10'sd491, 11'sd-932}, {12'sd1302, 11'sd516, 13'sd-3206}, {13'sd2398, 10'sd-294, 12'sd-1035}},
{{13'sd2815, 10'sd-400, 13'sd-2580}, {9'sd-135, 12'sd1811, 10'sd-472}, {13'sd2407, 13'sd-2713, 10'sd-467}},
{{12'sd1397, 12'sd-1825, 13'sd2109}, {12'sd-1389, 13'sd2106, 12'sd-2045}, {11'sd674, 13'sd-2221, 11'sd670}},
{{12'sd-1132, 8'sd-66, 11'sd-917}, {12'sd-1118, 13'sd-2733, 12'sd-1658}, {12'sd-1078, 12'sd1500, 11'sd-614}},
{{13'sd2589, 13'sd-2286, 11'sd791}, {12'sd-1426, 13'sd-2137, 11'sd802}, {12'sd-1359, 12'sd1100, 12'sd-1354}},
{{12'sd-1833, 13'sd-2639, 13'sd2341}, {12'sd1874, 10'sd-467, 12'sd1586}, {12'sd1333, 13'sd-2159, 13'sd-2330}},
{{9'sd156, 13'sd-2177, 11'sd-865}, {10'sd-332, 13'sd-2264, 13'sd-2103}, {12'sd-1584, 12'sd-1199, 12'sd-1989}},
{{10'sd303, 13'sd2262, 10'sd373}, {11'sd988, 12'sd-1939, 12'sd-1369}, {12'sd1578, 11'sd618, 12'sd-1142}},
{{13'sd3176, 11'sd-522, 13'sd2200}, {13'sd3085, 13'sd2147, 10'sd-335}, {12'sd1833, 9'sd-132, 12'sd-1368}},
{{13'sd-2246, 7'sd-34, 10'sd333}, {11'sd871, 11'sd-967, 11'sd852}, {11'sd-804, 12'sd-1671, 12'sd1728}},
{{14'sd-6164, 11'sd963, 12'sd-1218}, {13'sd-3727, 10'sd-458, 12'sd1506}, {13'sd-2951, 11'sd-1005, 12'sd1113}},
{{13'sd2103, 11'sd593, 13'sd2404}, {12'sd1932, 12'sd-1865, 9'sd130}, {11'sd901, 12'sd1183, 11'sd609}},
{{13'sd2282, 12'sd1044, 11'sd830}, {13'sd-2312, 12'sd-1473, 13'sd-2709}, {11'sd-563, 11'sd927, 8'sd-127}},
{{12'sd1916, 11'sd-546, 13'sd2657}, {12'sd1816, 11'sd-811, 10'sd-283}, {12'sd1553, 13'sd2104, 13'sd3210}},
{{12'sd1504, 12'sd-1573, 12'sd-1348}, {12'sd-1075, 13'sd2781, 12'sd-1506}, {12'sd-1123, 12'sd-1084, 13'sd2369}},
{{11'sd655, 12'sd-1477, 12'sd-1443}, {12'sd-1237, 13'sd-2987, 11'sd-923}, {11'sd756, 12'sd1641, 13'sd-2762}},
{{12'sd-1831, 11'sd-623, 13'sd-2589}, {11'sd846, 12'sd1295, 12'sd1643}, {13'sd-2536, 8'sd120, 9'sd191}},
{{13'sd2954, 12'sd1964, 12'sd-1918}, {12'sd-1845, 12'sd1678, 13'sd-2434}, {12'sd-1529, 14'sd-4703, 13'sd-2648}},
{{11'sd-667, 13'sd2071, 12'sd-1864}, {12'sd1100, 11'sd870, 5'sd-14}, {12'sd-1347, 12'sd1822, 10'sd-284}},
{{13'sd-2867, 11'sd-637, 12'sd1866}, {11'sd765, 11'sd746, 13'sd2090}, {11'sd-664, 12'sd-1792, 12'sd-1616}},
{{12'sd1822, 13'sd2497, 9'sd-219}, {12'sd1458, 10'sd498, 9'sd-213}, {11'sd-536, 11'sd-910, 13'sd2478}},
{{12'sd-1537, 10'sd330, 11'sd-974}, {12'sd-1887, 12'sd1894, 12'sd-1835}, {14'sd-4096, 11'sd-765, 12'sd-1165}},
{{13'sd2341, 13'sd2201, 12'sd-1979}, {12'sd-1411, 9'sd197, 11'sd811}, {8'sd125, 12'sd1847, 13'sd-2925}},
{{12'sd1750, 13'sd2736, 10'sd439}, {12'sd1866, 12'sd-1106, 11'sd692}, {12'sd-1973, 13'sd-2649, 13'sd2404}},
{{11'sd575, 12'sd-1620, 13'sd-2608}, {12'sd-1824, 12'sd-1265, 11'sd-824}, {14'sd4142, 13'sd2255, 13'sd2296}},
{{13'sd-2656, 10'sd429, 11'sd-925}, {13'sd-2347, 13'sd-2152, 11'sd761}, {12'sd-1857, 13'sd2406, 7'sd47}},
{{10'sd-270, 9'sd-138, 11'sd529}, {12'sd-1780, 12'sd1250, 12'sd-1988}, {12'sd1877, 12'sd-1246, 12'sd1414}},
{{12'sd2039, 13'sd2146, 9'sd201}, {11'sd-883, 13'sd-2049, 12'sd1491}, {12'sd1270, 8'sd-80, 10'sd489}},
{{11'sd843, 12'sd1498, 10'sd493}, {9'sd173, 11'sd828, 8'sd-64}, {13'sd-3444, 11'sd-608, 12'sd1810}},
{{13'sd-2691, 11'sd674, 13'sd3294}, {8'sd-71, 11'sd877, 11'sd606}, {12'sd-1715, 12'sd2011, 11'sd-592}},
{{12'sd1953, 11'sd-776, 11'sd-920}, {1'sd0, 12'sd1245, 5'sd11}, {12'sd-1567, 13'sd-2575, 13'sd2273}},
{{12'sd1571, 12'sd-2030, 12'sd-1417}, {12'sd-1074, 13'sd-2415, 13'sd-3546}, {13'sd2569, 12'sd1543, 13'sd-2464}},
{{13'sd-2330, 11'sd798, 12'sd-1314}, {12'sd-1930, 13'sd-2116, 11'sd-767}, {13'sd2123, 12'sd-1373, 11'sd-677}},
{{12'sd1797, 8'sd95, 12'sd-1182}, {12'sd-1602, 12'sd-1821, 12'sd-1466}, {13'sd-2137, 12'sd2046, 13'sd2386}},
{{11'sd-667, 13'sd2139, 11'sd-762}, {11'sd-926, 9'sd132, 11'sd-599}, {12'sd-1793, 13'sd2670, 13'sd2091}},
{{12'sd-1583, 13'sd2772, 13'sd2707}, {12'sd1736, 13'sd-2607, 13'sd2302}, {13'sd-2190, 7'sd57, 10'sd-348}},
{{11'sd-807, 12'sd1540, 13'sd2901}, {13'sd-2196, 13'sd2095, 10'sd435}, {13'sd-3487, 12'sd1827, 10'sd-320}},
{{13'sd4049, 12'sd-1222, 13'sd2136}, {11'sd-827, 12'sd1292, 12'sd-1582}, {12'sd2029, 9'sd-176, 11'sd874}},
{{12'sd-1632, 12'sd-1253, 12'sd1747}, {13'sd2156, 13'sd2207, 12'sd-1078}, {10'sd-361, 12'sd1252, 11'sd-955}},
{{11'sd612, 10'sd-450, 7'sd46}, {10'sd475, 12'sd1615, 12'sd-1096}, {12'sd1693, 12'sd-1033, 8'sd-107}},
{{13'sd2182, 12'sd1780, 12'sd1623}, {12'sd1969, 10'sd420, 13'sd-2117}, {10'sd261, 10'sd415, 13'sd-2218}},
{{12'sd1047, 10'sd440, 12'sd1100}, {12'sd-1532, 11'sd-628, 11'sd-724}, {11'sd887, 12'sd-1360, 12'sd-1839}},
{{11'sd-888, 12'sd-1049, 12'sd1497}, {10'sd473, 13'sd2688, 10'sd374}, {7'sd57, 11'sd691, 11'sd524}},
{{12'sd-1627, 10'sd323, 11'sd760}, {13'sd-2975, 12'sd1040, 12'sd1982}, {11'sd-724, 13'sd3498, 12'sd-1440}},
{{12'sd-1128, 8'sd77, 13'sd-2340}, {12'sd1477, 12'sd1317, 13'sd2533}, {12'sd1463, 10'sd268, 11'sd724}},
{{11'sd833, 10'sd-283, 12'sd-1330}, {13'sd-2129, 6'sd-29, 12'sd1631}, {12'sd-1840, 10'sd-470, 13'sd2678}},
{{12'sd-1373, 12'sd-1054, 13'sd-2497}, {12'sd-1077, 12'sd1854, 12'sd-1808}, {13'sd-2202, 13'sd-2123, 12'sd-1892}},
{{13'sd-2409, 12'sd1159, 13'sd2350}, {12'sd-1276, 11'sd706, 11'sd681}, {12'sd-1475, 11'sd707, 11'sd-769}},
{{13'sd2566, 13'sd2368, 10'sd396}, {12'sd1876, 7'sd-43, 8'sd69}, {13'sd2626, 9'sd173, 11'sd-643}},
{{12'sd-1337, 13'sd2887, 12'sd1517}, {11'sd-958, 12'sd-1201, 12'sd-1649}, {13'sd-2275, 8'sd122, 12'sd-1671}},
{{12'sd-1860, 12'sd-1262, 8'sd112}, {11'sd-930, 6'sd21, 11'sd625}, {11'sd841, 12'sd-1950, 13'sd2205}},
{{13'sd-2548, 11'sd-801, 13'sd2628}, {12'sd1652, 13'sd2141, 13'sd-2720}, {13'sd-2615, 12'sd-1674, 11'sd859}},
{{11'sd980, 11'sd-856, 13'sd2600}, {12'sd-1152, 12'sd-1353, 11'sd833}, {12'sd-1381, 12'sd-1718, 4'sd-7}},
{{10'sd385, 10'sd311, 11'sd1018}, {10'sd-261, 12'sd1920, 12'sd1912}, {12'sd1242, 13'sd-3017, 11'sd746}},
{{11'sd870, 12'sd-1189, 12'sd-1387}, {12'sd-1307, 11'sd-521, 12'sd-1267}, {12'sd1916, 13'sd-2071, 13'sd-2250}},
{{11'sd760, 12'sd1053, 12'sd-1871}, {13'sd2327, 11'sd-818, 13'sd-2239}, {13'sd2712, 12'sd-1148, 13'sd2059}},
{{13'sd2067, 10'sd-390, 11'sd969}, {11'sd-623, 12'sd1982, 11'sd-613}, {12'sd-1766, 12'sd1374, 12'sd1925}},
{{13'sd3791, 11'sd-631, 13'sd2538}, {13'sd3742, 10'sd-316, 12'sd1616}, {14'sd4332, 11'sd-601, 8'sd-95}},
{{13'sd-2302, 10'sd-308, 11'sd-789}, {11'sd758, 13'sd-2513, 11'sd811}, {12'sd1811, 12'sd-1961, 13'sd2184}},
{{10'sd452, 13'sd-2377, 13'sd2522}, {9'sd139, 11'sd870, 11'sd-638}, {12'sd1784, 12'sd-1237, 12'sd1824}},
{{12'sd-1095, 12'sd1621, 12'sd-2012}, {8'sd-79, 13'sd-2479, 12'sd1740}, {11'sd664, 12'sd1232, 9'sd-137}},
{{12'sd-1376, 13'sd-2179, 12'sd-1843}, {12'sd-1180, 13'sd-2188, 13'sd-2069}, {8'sd72, 13'sd2408, 8'sd89}},
{{12'sd-1773, 10'sd404, 12'sd1245}, {13'sd-2992, 12'sd-1501, 10'sd289}, {13'sd2456, 12'sd1846, 13'sd-2498}},
{{4'sd-4, 12'sd-1502, 11'sd637}, {12'sd1336, 12'sd-1885, 13'sd2357}, {11'sd-547, 13'sd-2563, 6'sd19}}},
{
{{12'sd-1865, 11'sd609, 13'sd-2086}, {12'sd-1938, 13'sd2381, 12'sd-1447}, {13'sd-2544, 11'sd-629, 12'sd-1632}},
{{13'sd-2726, 8'sd65, 12'sd1377}, {9'sd-142, 12'sd-1515, 12'sd-1593}, {13'sd-2882, 13'sd-2485, 13'sd-2879}},
{{11'sd937, 9'sd-165, 11'sd980}, {11'sd-737, 13'sd-3294, 12'sd1922}, {12'sd-1091, 11'sd973, 6'sd23}},
{{11'sd1020, 10'sd-293, 12'sd-2042}, {13'sd2425, 12'sd-1729, 13'sd2524}, {11'sd-794, 12'sd1159, 13'sd2462}},
{{13'sd-2808, 13'sd2373, 12'sd1889}, {13'sd-2089, 13'sd-2175, 12'sd-1645}, {10'sd-430, 12'sd1210, 13'sd-2203}},
{{12'sd1269, 10'sd509, 12'sd2003}, {9'sd165, 12'sd-1245, 13'sd2281}, {11'sd-723, 12'sd1471, 13'sd2573}},
{{13'sd2434, 12'sd1576, 12'sd1154}, {12'sd-1325, 12'sd-1455, 11'sd-629}, {13'sd-2451, 12'sd1910, 12'sd1549}},
{{12'sd1364, 12'sd-1991, 12'sd1965}, {7'sd-53, 8'sd101, 12'sd1378}, {12'sd-2029, 10'sd383, 12'sd1747}},
{{12'sd-1902, 11'sd-1021, 11'sd756}, {12'sd-1946, 12'sd-1276, 13'sd-2466}, {12'sd1661, 11'sd-602, 12'sd-1366}},
{{13'sd2361, 11'sd576, 12'sd1303}, {13'sd-2225, 12'sd-1676, 13'sd-2666}, {12'sd-1390, 11'sd-757, 11'sd640}},
{{12'sd-1831, 11'sd-799, 10'sd266}, {12'sd1051, 12'sd1182, 8'sd99}, {9'sd-169, 11'sd627, 11'sd-599}},
{{11'sd-917, 11'sd-563, 12'sd-1967}, {9'sd-184, 12'sd1033, 11'sd833}, {7'sd-32, 10'sd458, 12'sd1947}},
{{11'sd-664, 9'sd213, 8'sd-120}, {12'sd1587, 13'sd-2089, 13'sd-2602}, {9'sd-149, 12'sd-1448, 9'sd203}},
{{11'sd748, 13'sd2097, 8'sd83}, {12'sd1639, 12'sd-1059, 11'sd-932}, {13'sd-2477, 12'sd-1716, 11'sd970}},
{{12'sd1581, 12'sd-1876, 13'sd-2673}, {12'sd-1102, 10'sd365, 11'sd-656}, {12'sd1403, 11'sd782, 12'sd-1882}},
{{13'sd-2629, 12'sd1075, 11'sd882}, {11'sd-896, 12'sd1768, 12'sd-1220}, {12'sd1520, 12'sd1933, 11'sd-531}},
{{13'sd-2874, 11'sd-607, 12'sd-1763}, {12'sd-1812, 9'sd-244, 12'sd1375}, {7'sd53, 12'sd1820, 13'sd3436}},
{{11'sd568, 12'sd-1139, 13'sd2416}, {12'sd1190, 13'sd-3615, 9'sd174}, {12'sd-1643, 13'sd-2244, 11'sd873}},
{{11'sd536, 12'sd-1408, 5'sd-9}, {11'sd-839, 10'sd472, 9'sd159}, {9'sd-180, 9'sd-238, 7'sd61}},
{{11'sd712, 9'sd223, 9'sd240}, {11'sd550, 10'sd-373, 12'sd-1830}, {13'sd2732, 13'sd3594, 10'sd330}},
{{13'sd-2589, 9'sd220, 12'sd1629}, {12'sd-1223, 10'sd-339, 12'sd-1407}, {10'sd361, 13'sd2230, 11'sd-700}},
{{12'sd-1176, 13'sd-2166, 11'sd567}, {8'sd103, 7'sd-34, 12'sd1439}, {13'sd-2505, 12'sd-1306, 9'sd-146}},
{{13'sd2106, 11'sd-988, 12'sd1123}, {12'sd-1702, 12'sd-1835, 11'sd-704}, {11'sd-712, 11'sd714, 11'sd-730}},
{{10'sd465, 12'sd-1925, 12'sd-1511}, {13'sd-2506, 12'sd1691, 12'sd1164}, {12'sd-1952, 11'sd543, 13'sd-2172}},
{{11'sd-858, 11'sd1006, 13'sd2406}, {13'sd2959, 10'sd469, 13'sd-2511}, {8'sd111, 14'sd-4156, 12'sd-1475}},
{{10'sd410, 11'sd-895, 12'sd1250}, {8'sd-107, 12'sd-1133, 12'sd-1247}, {13'sd2663, 13'sd2359, 11'sd-863}},
{{13'sd2503, 13'sd2211, 13'sd-2394}, {8'sd124, 13'sd2649, 12'sd2028}, {13'sd-2395, 12'sd-1953, 13'sd-2395}},
{{13'sd2423, 12'sd-1375, 12'sd-1704}, {12'sd-1310, 13'sd-2129, 11'sd987}, {13'sd2454, 9'sd200, 11'sd673}},
{{13'sd2301, 13'sd-2106, 11'sd-631}, {13'sd-2718, 10'sd-411, 10'sd487}, {13'sd2429, 13'sd2622, 11'sd892}},
{{13'sd-2687, 11'sd-718, 11'sd-916}, {12'sd-1215, 12'sd1289, 12'sd-1552}, {9'sd144, 13'sd2600, 13'sd3314}},
{{12'sd1842, 12'sd1691, 8'sd-80}, {12'sd1283, 13'sd2426, 11'sd-843}, {13'sd2609, 12'sd-1610, 12'sd-1567}},
{{12'sd1550, 11'sd1013, 12'sd-1285}, {12'sd1424, 12'sd-1440, 13'sd-2780}, {12'sd-1166, 11'sd688, 11'sd918}},
{{13'sd2365, 13'sd-2885, 13'sd2364}, {12'sd1985, 12'sd1025, 13'sd-2484}, {13'sd-2148, 10'sd-364, 12'sd-1338}},
{{11'sd559, 13'sd-2356, 12'sd1545}, {13'sd3039, 13'sd-2416, 9'sd201}, {11'sd-682, 11'sd779, 12'sd1608}},
{{11'sd-880, 12'sd1158, 13'sd2558}, {10'sd492, 11'sd-738, 12'sd1973}, {12'sd1078, 11'sd-637, 12'sd-1720}},
{{13'sd2152, 11'sd764, 13'sd-2138}, {11'sd755, 5'sd13, 13'sd2454}, {11'sd-662, 13'sd-2214, 12'sd-1456}},
{{13'sd-2426, 12'sd1514, 12'sd-1568}, {12'sd1864, 12'sd1647, 10'sd-398}, {10'sd448, 9'sd233, 12'sd1878}},
{{13'sd-4022, 10'sd-435, 11'sd611}, {13'sd-2054, 10'sd-285, 13'sd-2512}, {13'sd-3922, 12'sd-1636, 12'sd1984}},
{{11'sd-959, 13'sd-2539, 12'sd1649}, {10'sd473, 12'sd1291, 11'sd1006}, {12'sd-1569, 13'sd2847, 13'sd2658}},
{{10'sd449, 13'sd2460, 12'sd1383}, {11'sd-619, 12'sd-1159, 11'sd-936}, {12'sd1330, 13'sd-2059, 13'sd-2135}},
{{11'sd895, 12'sd-1206, 11'sd-615}, {11'sd-828, 9'sd-187, 11'sd805}, {10'sd425, 13'sd-2601, 8'sd71}},
{{11'sd-704, 13'sd2530, 13'sd2859}, {13'sd-2390, 9'sd228, 13'sd-2390}, {12'sd-1746, 12'sd-1705, 11'sd-1010}},
{{9'sd-129, 12'sd-1954, 12'sd1804}, {13'sd-2796, 12'sd-1289, 13'sd-2169}, {11'sd-629, 12'sd-1627, 12'sd1270}},
{{12'sd-1538, 13'sd3221, 11'sd970}, {13'sd2593, 13'sd3468, 13'sd2237}, {12'sd-1373, 13'sd3336, 13'sd2945}},
{{11'sd809, 13'sd-2482, 3'sd-2}, {12'sd1473, 11'sd568, 12'sd-1722}, {10'sd327, 12'sd-1334, 11'sd-683}},
{{12'sd-1658, 13'sd-2880, 13'sd-2514}, {12'sd1935, 9'sd-245, 10'sd295}, {12'sd1208, 13'sd-3001, 12'sd-1609}},
{{10'sd-274, 13'sd2291, 13'sd-2078}, {9'sd-214, 13'sd-2104, 12'sd1377}, {13'sd-2134, 11'sd935, 12'sd1726}},
{{12'sd-1983, 12'sd1919, 12'sd1631}, {12'sd-1355, 12'sd1222, 11'sd-963}, {12'sd1278, 12'sd-1366, 12'sd-1913}},
{{12'sd-1980, 12'sd-1148, 12'sd-1347}, {12'sd1708, 12'sd-2046, 12'sd-1553}, {11'sd632, 12'sd-1565, 13'sd-2104}},
{{12'sd2044, 12'sd-1572, 11'sd697}, {11'sd-811, 2'sd1, 12'sd-1612}, {12'sd1363, 13'sd-2168, 13'sd2521}},
{{13'sd-2577, 12'sd-1501, 10'sd447}, {13'sd-2341, 13'sd-2358, 12'sd1388}, {12'sd-1528, 12'sd-1060, 10'sd283}},
{{12'sd1426, 12'sd-1483, 12'sd-1254}, {13'sd2709, 7'sd46, 12'sd-1039}, {12'sd1899, 10'sd-267, 11'sd-837}},
{{11'sd563, 9'sd128, 13'sd2598}, {13'sd-2896, 11'sd-576, 12'sd-1667}, {13'sd-3469, 13'sd-3112, 12'sd1525}},
{{8'sd-100, 13'sd2827, 12'sd-1880}, {13'sd2895, 12'sd-1419, 11'sd932}, {12'sd1748, 11'sd527, 12'sd1482}},
{{13'sd-2086, 12'sd1999, 12'sd-1558}, {13'sd2887, 12'sd-1252, 12'sd1621}, {13'sd2053, 13'sd-2062, 13'sd2373}},
{{12'sd1886, 9'sd-212, 13'sd2100}, {12'sd1106, 12'sd1832, 9'sd-245}, {9'sd141, 13'sd2654, 12'sd-1576}},
{{13'sd-2078, 12'sd-1996, 12'sd1410}, {12'sd-1608, 12'sd1182, 11'sd682}, {12'sd1783, 13'sd-2177, 13'sd-2456}},
{{12'sd1143, 13'sd2326, 11'sd564}, {12'sd-1585, 9'sd176, 12'sd-2044}, {13'sd-2572, 11'sd-886, 10'sd-457}},
{{13'sd2811, 11'sd1021, 12'sd-1856}, {13'sd2348, 12'sd-1715, 8'sd119}, {13'sd2240, 11'sd790, 12'sd-1058}},
{{11'sd-554, 12'sd-2034, 12'sd1560}, {13'sd-2235, 13'sd-2684, 12'sd1934}, {12'sd-1368, 12'sd1545, 13'sd-2138}},
{{11'sd-871, 12'sd1182, 11'sd-777}, {13'sd2653, 13'sd-2078, 11'sd-614}, {13'sd2769, 12'sd1750, 12'sd1835}},
{{11'sd-651, 10'sd-507, 11'sd-706}, {12'sd1169, 9'sd-228, 12'sd1905}, {13'sd-2289, 11'sd-697, 13'sd2915}},
{{11'sd760, 13'sd2144, 11'sd721}, {12'sd-1024, 11'sd-810, 12'sd-1094}, {10'sd310, 12'sd-2043, 10'sd328}},
{{12'sd2005, 13'sd-2064, 9'sd254}, {13'sd2223, 12'sd-1816, 13'sd2126}, {10'sd-425, 13'sd-2344, 13'sd2963}}},
{
{{12'sd-1716, 10'sd-334, 11'sd-946}, {12'sd-1198, 11'sd734, 12'sd-1796}, {13'sd3195, 9'sd178, 13'sd2529}},
{{10'sd473, 12'sd-1752, 12'sd-1429}, {12'sd-1438, 9'sd176, 10'sd-266}, {12'sd-1293, 13'sd2133, 12'sd-1832}},
{{12'sd-1745, 8'sd-98, 12'sd-1986}, {12'sd1265, 13'sd2344, 11'sd634}, {12'sd-1289, 12'sd1412, 12'sd-1813}},
{{13'sd-2663, 12'sd-1850, 13'sd-2096}, {13'sd2106, 13'sd2430, 13'sd2474}, {11'sd963, 12'sd1230, 10'sd380}},
{{11'sd750, 11'sd521, 12'sd1281}, {13'sd-2529, 11'sd558, 13'sd-2511}, {12'sd1811, 13'sd3660, 11'sd-643}},
{{12'sd1822, 13'sd-2194, 11'sd-535}, {11'sd910, 10'sd-453, 12'sd1540}, {12'sd1507, 13'sd-2463, 9'sd161}},
{{13'sd-3646, 13'sd-3232, 12'sd-1650}, {12'sd-1491, 12'sd-1579, 13'sd-2663}, {13'sd-2300, 12'sd1337, 12'sd-1244}},
{{12'sd-1358, 11'sd-653, 8'sd-126}, {13'sd-2883, 8'sd123, 10'sd437}, {12'sd1227, 13'sd3561, 11'sd-587}},
{{11'sd537, 12'sd1429, 13'sd2953}, {13'sd2471, 12'sd-1857, 13'sd2542}, {13'sd3720, 12'sd1427, 13'sd2799}},
{{12'sd-1361, 10'sd-377, 11'sd-938}, {13'sd-2361, 11'sd-877, 11'sd-527}, {13'sd-2672, 12'sd-1415, 11'sd769}},
{{12'sd1561, 9'sd-246, 11'sd-761}, {12'sd1128, 12'sd1037, 12'sd-1524}, {14'sd-4524, 12'sd-1563, 12'sd-1589}},
{{10'sd464, 13'sd-2455, 12'sd-1375}, {10'sd-346, 13'sd2324, 10'sd257}, {12'sd1825, 9'sd236, 12'sd1797}},
{{10'sd-266, 11'sd-842, 10'sd-487}, {12'sd1118, 11'sd-903, 8'sd-71}, {12'sd-1994, 11'sd-898, 12'sd1510}},
{{12'sd-1327, 12'sd-1275, 12'sd-1516}, {10'sd316, 12'sd1491, 12'sd1068}, {12'sd-1677, 13'sd-2544, 13'sd-2336}},
{{13'sd2836, 11'sd-970, 11'sd1016}, {12'sd1041, 11'sd877, 9'sd-241}, {13'sd-2348, 12'sd-1671, 12'sd1438}},
{{11'sd-554, 12'sd-1777, 12'sd1706}, {13'sd-2971, 12'sd-1033, 12'sd-1058}, {13'sd2465, 12'sd1766, 13'sd2952}},
{{12'sd-1636, 8'sd116, 13'sd-2890}, {11'sd-678, 10'sd397, 11'sd-874}, {12'sd-1968, 12'sd1898, 12'sd-2032}},
{{14'sd-5474, 8'sd-119, 13'sd-3403}, {13'sd-2528, 12'sd1417, 10'sd279}, {13'sd-2180, 10'sd396, 13'sd3087}},
{{12'sd-1491, 12'sd-1439, 11'sd947}, {13'sd-2334, 13'sd2203, 11'sd897}, {11'sd663, 12'sd1141, 7'sd-48}},
{{13'sd-2225, 13'sd-2224, 12'sd1620}, {12'sd-1612, 12'sd-1411, 12'sd-1407}, {13'sd-2915, 12'sd-1531, 12'sd1193}},
{{13'sd2472, 13'sd2689, 12'sd-1246}, {12'sd1330, 11'sd854, 13'sd-2410}, {12'sd2020, 11'sd-693, 12'sd-2026}},
{{12'sd1873, 10'sd393, 13'sd2062}, {10'sd306, 12'sd1738, 13'sd2260}, {8'sd-68, 10'sd446, 12'sd-1503}},
{{10'sd-450, 11'sd-1009, 11'sd801}, {12'sd1097, 13'sd2258, 13'sd-2124}, {10'sd350, 13'sd-2686, 12'sd1979}},
{{9'sd-138, 10'sd-467, 12'sd-1066}, {12'sd-1992, 10'sd-421, 13'sd-2439}, {11'sd-999, 8'sd-95, 12'sd1464}},
{{11'sd944, 13'sd2659, 13'sd2591}, {14'sd4168, 13'sd2834, 12'sd1770}, {13'sd3004, 11'sd-679, 12'sd1188}},
{{12'sd1685, 12'sd-1966, 13'sd2448}, {13'sd-2567, 12'sd1675, 7'sd-32}, {12'sd1811, 12'sd-1554, 13'sd2484}},
{{9'sd-218, 10'sd-401, 12'sd1674}, {9'sd139, 8'sd-109, 10'sd329}, {12'sd1992, 12'sd1621, 11'sd850}},
{{12'sd-1811, 12'sd-1912, 13'sd2611}, {10'sd-355, 12'sd-1068, 12'sd1402}, {12'sd1850, 10'sd461, 12'sd-1484}},
{{13'sd-2590, 10'sd-359, 12'sd-1948}, {12'sd-1440, 11'sd-1002, 10'sd497}, {13'sd-3160, 12'sd1993, 12'sd-1567}},
{{12'sd-1185, 12'sd-1404, 12'sd1255}, {12'sd1263, 13'sd2141, 13'sd2854}, {10'sd291, 12'sd-1848, 9'sd136}},
{{12'sd1549, 12'sd1622, 12'sd1568}, {12'sd-1885, 13'sd-2053, 7'sd33}, {12'sd1447, 12'sd1873, 12'sd-2009}},
{{12'sd-1708, 11'sd-538, 13'sd-3490}, {12'sd1049, 12'sd1405, 13'sd-2141}, {13'sd3610, 13'sd2484, 12'sd-1866}},
{{12'sd1367, 9'sd179, 12'sd-1275}, {10'sd-385, 11'sd882, 11'sd870}, {11'sd-623, 9'sd245, 11'sd-985}},
{{12'sd-1863, 11'sd598, 12'sd-1855}, {11'sd-753, 7'sd61, 12'sd1560}, {11'sd-863, 13'sd-3252, 11'sd-728}},
{{12'sd-1097, 8'sd-102, 12'sd-1640}, {11'sd-715, 10'sd-485, 12'sd-1462}, {13'sd2393, 10'sd310, 13'sd2469}},
{{12'sd-1257, 12'sd-1513, 11'sd631}, {9'sd211, 13'sd2277, 8'sd112}, {13'sd2223, 13'sd-2436, 12'sd1426}},
{{11'sd-545, 11'sd606, 13'sd-2390}, {10'sd328, 13'sd-2147, 7'sd39}, {12'sd1627, 9'sd-144, 13'sd2129}},
{{12'sd-1843, 9'sd-254, 12'sd-1184}, {11'sd-886, 14'sd4295, 11'sd-777}, {13'sd2075, 14'sd4713, 11'sd774}},
{{12'sd1159, 13'sd-2474, 14'sd-4764}, {10'sd-303, 12'sd-1263, 13'sd-2388}, {10'sd-356, 13'sd2324, 12'sd1500}},
{{13'sd-3277, 12'sd-2023, 12'sd-1342}, {12'sd-1498, 11'sd-691, 12'sd-1051}, {12'sd-1237, 13'sd2988, 13'sd2891}},
{{13'sd2310, 13'sd-2447, 11'sd-571}, {13'sd-2111, 11'sd-670, 12'sd-1054}, {12'sd-1152, 8'sd80, 13'sd-2064}},
{{10'sd448, 13'sd-2365, 11'sd-964}, {6'sd28, 11'sd-933, 13'sd-2212}, {12'sd-1458, 13'sd2442, 12'sd1046}},
{{11'sd-720, 13'sd-2748, 12'sd1150}, {10'sd320, 10'sd485, 12'sd-1271}, {12'sd-1791, 9'sd-171, 13'sd2056}},
{{13'sd3124, 11'sd-631, 13'sd2261}, {13'sd2704, 12'sd1320, 13'sd2945}, {9'sd190, 7'sd42, 8'sd91}},
{{12'sd-1627, 11'sd550, 13'sd2124}, {13'sd-2117, 12'sd-1134, 13'sd2857}, {12'sd-1371, 12'sd-1217, 12'sd-1100}},
{{12'sd1760, 13'sd2307, 13'sd2343}, {11'sd783, 12'sd1299, 12'sd-1573}, {12'sd1661, 12'sd-1457, 9'sd220}},
{{12'sd-1432, 11'sd-632, 13'sd-2349}, {11'sd927, 13'sd3161, 10'sd-303}, {12'sd-1081, 12'sd1774, 12'sd-1859}},
{{12'sd1476, 12'sd-1894, 10'sd-306}, {10'sd-492, 12'sd1169, 13'sd-2140}, {11'sd-965, 13'sd-2398, 12'sd-1716}},
{{12'sd-1881, 13'sd2103, 11'sd-527}, {13'sd-2450, 10'sd-328, 11'sd-992}, {10'sd-371, 12'sd-1446, 12'sd1826}},
{{11'sd-645, 12'sd-1117, 7'sd53}, {10'sd-435, 9'sd235, 11'sd-629}, {12'sd-1121, 10'sd303, 13'sd-2353}},
{{11'sd-568, 12'sd1490, 12'sd-1818}, {10'sd-320, 12'sd1466, 13'sd2454}, {13'sd2175, 12'sd-1493, 13'sd-2652}},
{{12'sd-1125, 12'sd-1419, 13'sd2515}, {8'sd-95, 12'sd-1689, 11'sd-908}, {12'sd-1978, 11'sd-840, 9'sd181}},
{{11'sd887, 13'sd-3006, 13'sd-3983}, {13'sd3157, 11'sd-825, 8'sd112}, {11'sd910, 13'sd3847, 9'sd-129}},
{{8'sd79, 13'sd2387, 12'sd-1229}, {11'sd625, 13'sd2757, 12'sd1935}, {12'sd1753, 13'sd2233, 12'sd1959}},
{{12'sd-1921, 12'sd1026, 5'sd-13}, {10'sd288, 13'sd-2316, 11'sd746}, {12'sd1263, 12'sd1314, 11'sd-810}},
{{12'sd1928, 12'sd-1137, 10'sd-287}, {13'sd2401, 13'sd-2140, 13'sd-2537}, {13'sd-2119, 12'sd1467, 13'sd-2366}},
{{12'sd1388, 11'sd-645, 11'sd-986}, {11'sd-701, 12'sd1223, 12'sd-2045}, {13'sd2141, 10'sd500, 10'sd-481}},
{{10'sd-449, 10'sd277, 12'sd-1825}, {11'sd948, 12'sd-1316, 12'sd1434}, {14'sd4772, 13'sd-2278, 12'sd1287}},
{{11'sd542, 13'sd3366, 12'sd1734}, {13'sd2828, 13'sd3603, 9'sd-253}, {11'sd945, 8'sd116, 12'sd-1175}},
{{12'sd-1988, 11'sd-793, 13'sd2448}, {12'sd-1076, 11'sd-801, 11'sd-851}, {10'sd-453, 12'sd-1757, 13'sd2907}},
{{12'sd-1635, 8'sd117, 13'sd-2049}, {12'sd-1162, 13'sd2665, 11'sd723}, {13'sd3082, 13'sd3465, 11'sd-840}},
{{11'sd-1018, 13'sd-2368, 7'sd57}, {13'sd-2540, 12'sd1127, 12'sd-1822}, {13'sd2317, 13'sd-2093, 13'sd-2355}},
{{11'sd528, 12'sd1876, 8'sd-68}, {12'sd-1891, 12'sd1178, 13'sd-2876}, {13'sd2478, 12'sd1553, 13'sd-2304}},
{{12'sd-1713, 13'sd2201, 11'sd805}, {13'sd2051, 13'sd3351, 12'sd1535}, {13'sd2736, 12'sd1480, 13'sd2430}}},
{
{{12'sd-1632, 13'sd-2831, 13'sd-3316}, {12'sd1050, 13'sd-3473, 13'sd-2878}, {10'sd423, 9'sd-222, 13'sd-3159}},
{{12'sd-1655, 11'sd-617, 13'sd2135}, {12'sd1547, 10'sd387, 12'sd-1923}, {13'sd-2622, 13'sd-2914, 10'sd394}},
{{10'sd-428, 12'sd-1678, 10'sd287}, {13'sd2329, 10'sd-343, 13'sd3590}, {13'sd2593, 13'sd2670, 13'sd2882}},
{{12'sd-1521, 11'sd-808, 13'sd-2160}, {12'sd1846, 13'sd2084, 12'sd-1577}, {12'sd1795, 12'sd1631, 13'sd-2867}},
{{12'sd1269, 11'sd1014, 10'sd-477}, {12'sd-1732, 12'sd1048, 11'sd916}, {13'sd2120, 12'sd1695, 12'sd1675}},
{{10'sd411, 11'sd879, 11'sd971}, {13'sd-2068, 10'sd301, 12'sd1889}, {13'sd2191, 13'sd2131, 9'sd172}},
{{13'sd3768, 9'sd-176, 10'sd427}, {12'sd-1824, 12'sd-1273, 13'sd2631}, {10'sd331, 12'sd1711, 12'sd-1631}},
{{13'sd2406, 11'sd978, 12'sd-1904}, {11'sd654, 13'sd-2307, 9'sd254}, {13'sd-2367, 13'sd-2209, 12'sd-2043}},
{{13'sd-2653, 7'sd57, 12'sd-1557}, {7'sd59, 11'sd541, 13'sd2259}, {8'sd91, 9'sd-235, 12'sd-1143}},
{{12'sd-1817, 12'sd1949, 13'sd2310}, {13'sd-2637, 12'sd-1814, 12'sd2019}, {11'sd-868, 13'sd-3088, 13'sd2210}},
{{13'sd2718, 13'sd2317, 13'sd-2545}, {13'sd2225, 12'sd2034, 13'sd-4057}, {12'sd1293, 12'sd-1266, 12'sd-2019}},
{{12'sd1583, 12'sd-1835, 13'sd-2209}, {12'sd1969, 8'sd-78, 12'sd-1888}, {12'sd2011, 13'sd2290, 13'sd-2460}},
{{11'sd665, 13'sd-2284, 14'sd4361}, {12'sd-1119, 12'sd-1924, 13'sd3321}, {9'sd-239, 10'sd357, 6'sd-25}},
{{13'sd2244, 13'sd2477, 12'sd1743}, {10'sd-341, 9'sd183, 11'sd1014}, {13'sd-2345, 8'sd-65, 12'sd-1454}},
{{9'sd-140, 13'sd2844, 11'sd570}, {11'sd-696, 13'sd2819, 12'sd-1355}, {11'sd-962, 12'sd1113, 12'sd1826}},
{{13'sd2828, 13'sd-2163, 13'sd-2450}, {13'sd2219, 13'sd2529, 12'sd1670}, {13'sd-2878, 13'sd-2483, 13'sd-2877}},
{{12'sd1626, 10'sd-425, 13'sd3634}, {12'sd1821, 12'sd1580, 12'sd-1507}, {7'sd36, 12'sd-1481, 10'sd353}},
{{12'sd-1831, 13'sd-3167, 9'sd-174}, {11'sd981, 12'sd-1797, 13'sd3930}, {14'sd4517, 12'sd1704, 13'sd2502}},
{{11'sd687, 12'sd-1780, 11'sd788}, {13'sd2335, 11'sd752, 12'sd-1545}, {11'sd-700, 11'sd-738, 12'sd1583}},
{{12'sd-1309, 13'sd2222, 12'sd1868}, {12'sd-1948, 12'sd-1660, 10'sd-260}, {13'sd-3323, 12'sd-1702, 13'sd-2238}},
{{11'sd578, 10'sd-384, 12'sd1984}, {11'sd554, 9'sd-187, 12'sd-1766}, {13'sd3063, 12'sd-1280, 13'sd3279}},
{{13'sd-2971, 10'sd311, 10'sd-277}, {13'sd-2590, 13'sd-2135, 12'sd1725}, {12'sd-1971, 12'sd-1556, 10'sd-498}},
{{12'sd-1486, 12'sd-1076, 13'sd-2313}, {12'sd1985, 11'sd598, 6'sd17}, {12'sd-1730, 13'sd2508, 11'sd942}},
{{12'sd-1173, 13'sd2062, 13'sd2324}, {12'sd-1795, 9'sd236, 12'sd-2014}, {12'sd1215, 13'sd2603, 11'sd646}},
{{13'sd-3500, 13'sd-2764, 12'sd1931}, {12'sd-2008, 12'sd-1467, 12'sd1818}, {14'sd4598, 12'sd1668, 14'sd4768}},
{{11'sd-584, 13'sd2769, 11'sd-643}, {10'sd498, 12'sd1156, 12'sd1070}, {11'sd-727, 12'sd1217, 11'sd-841}},
{{13'sd-2286, 13'sd2783, 13'sd-2944}, {12'sd1299, 13'sd2073, 12'sd-1570}, {10'sd-356, 12'sd-1338, 4'sd-6}},
{{10'sd414, 13'sd2075, 13'sd-2643}, {12'sd1324, 11'sd720, 10'sd456}, {10'sd274, 12'sd1835, 12'sd1465}},
{{11'sd-792, 13'sd2302, 11'sd-720}, {10'sd-468, 12'sd1096, 11'sd586}, {12'sd-1975, 11'sd-741, 11'sd666}},
{{12'sd-1844, 12'sd1338, 12'sd-1825}, {11'sd880, 12'sd1458, 6'sd31}, {13'sd-2228, 12'sd-1637, 11'sd886}},
{{13'sd-2249, 13'sd2208, 12'sd-1997}, {11'sd959, 8'sd85, 9'sd169}, {5'sd-13, 13'sd-2657, 11'sd958}},
{{10'sd355, 11'sd832, 13'sd-2730}, {10'sd310, 13'sd-3525, 13'sd-3467}, {12'sd-1649, 12'sd-1575, 12'sd-1234}},
{{13'sd-2870, 13'sd-2742, 12'sd-1902}, {9'sd174, 12'sd-1088, 11'sd-971}, {12'sd1920, 12'sd1450, 12'sd-2032}},
{{12'sd1028, 5'sd10, 12'sd2037}, {10'sd-352, 12'sd1348, 11'sd681}, {13'sd-2384, 12'sd1303, 12'sd-1747}},
{{11'sd-980, 11'sd-939, 13'sd-2487}, {10'sd509, 12'sd-1980, 12'sd1281}, {10'sd-511, 11'sd880, 12'sd-1819}},
{{12'sd1153, 12'sd-1121, 12'sd-1154}, {10'sd-383, 12'sd-1572, 8'sd115}, {12'sd1100, 13'sd2562, 11'sd940}},
{{12'sd1871, 11'sd635, 13'sd-2072}, {13'sd2638, 13'sd-2200, 12'sd-1569}, {13'sd3069, 11'sd-924, 13'sd2148}},
{{8'sd77, 12'sd1291, 13'sd-2544}, {12'sd1594, 12'sd1178, 13'sd-3915}, {11'sd825, 12'sd-1510, 13'sd-2779}},
{{13'sd2396, 12'sd-1315, 12'sd1874}, {12'sd-1401, 13'sd-3117, 12'sd-1399}, {13'sd-2352, 13'sd-2908, 12'sd1465}},
{{12'sd-1417, 13'sd-2295, 13'sd-2722}, {13'sd2948, 12'sd1056, 12'sd1063}, {13'sd2712, 12'sd1376, 10'sd499}},
{{13'sd3023, 7'sd-37, 11'sd-1015}, {11'sd512, 8'sd108, 12'sd-1955}, {11'sd638, 12'sd1287, 11'sd-891}},
{{13'sd-2138, 7'sd63, 11'sd-781}, {11'sd-948, 12'sd1876, 13'sd-2356}, {13'sd2290, 13'sd-2589, 12'sd-1287}},
{{13'sd2413, 11'sd749, 12'sd-1980}, {12'sd-1326, 12'sd1360, 13'sd-2168}, {12'sd-1817, 13'sd-2349, 13'sd-2144}},
{{12'sd-1683, 10'sd328, 12'sd-1288}, {12'sd1950, 13'sd2202, 13'sd-2396}, {13'sd-2645, 12'sd1893, 12'sd-1306}},
{{12'sd1250, 12'sd-1364, 12'sd1030}, {11'sd-831, 12'sd1556, 11'sd847}, {13'sd2519, 11'sd-812, 9'sd151}},
{{13'sd2048, 13'sd-2201, 10'sd-322}, {12'sd-1197, 11'sd698, 10'sd-403}, {9'sd-235, 13'sd2856, 10'sd321}},
{{12'sd1700, 13'sd2472, 13'sd2945}, {12'sd1565, 13'sd-2972, 10'sd-357}, {11'sd696, 13'sd2485, 13'sd2168}},
{{12'sd-1657, 11'sd-922, 12'sd1995}, {12'sd-1159, 11'sd-712, 10'sd-288}, {13'sd-2364, 13'sd2304, 12'sd1542}},
{{11'sd671, 11'sd-895, 11'sd756}, {8'sd-68, 11'sd991, 13'sd2088}, {10'sd-484, 9'sd-180, 13'sd-2531}},
{{7'sd41, 11'sd-572, 13'sd2695}, {12'sd-1840, 12'sd1266, 12'sd-1727}, {8'sd-127, 9'sd242, 13'sd2560}},
{{12'sd1509, 12'sd1225, 12'sd-1606}, {12'sd-1977, 12'sd2016, 12'sd1562}, {12'sd1173, 11'sd822, 10'sd-456}},
{{11'sd810, 10'sd-288, 12'sd1796}, {12'sd1854, 10'sd427, 12'sd1735}, {7'sd-40, 9'sd131, 12'sd-1912}},
{{12'sd1340, 11'sd967, 12'sd-1811}, {10'sd-411, 8'sd77, 9'sd-241}, {11'sd883, 13'sd4076, 13'sd3508}},
{{12'sd1908, 13'sd-3091, 11'sd-910}, {10'sd288, 12'sd1040, 13'sd-2284}, {12'sd1554, 12'sd-2035, 12'sd-1671}},
{{11'sd749, 13'sd2200, 12'sd1200}, {12'sd1429, 12'sd-1731, 11'sd822}, {12'sd-1206, 12'sd-1365, 12'sd1269}},
{{5'sd-15, 11'sd-570, 12'sd1144}, {12'sd1399, 13'sd2582, 13'sd-2427}, {13'sd2638, 12'sd-1518, 12'sd-1668}},
{{11'sd-533, 9'sd249, 12'sd-1082}, {12'sd1111, 12'sd-1183, 11'sd537}, {11'sd852, 12'sd1556, 13'sd3066}},
{{13'sd3157, 8'sd92, 11'sd-919}, {12'sd1357, 13'sd-3300, 13'sd-2235}, {14'sd5298, 12'sd2044, 12'sd1929}},
{{11'sd-860, 13'sd-3760, 13'sd-2413}, {11'sd572, 11'sd-714, 12'sd-1439}, {13'sd2458, 11'sd985, 12'sd-1074}},
{{12'sd1635, 12'sd1549, 11'sd-780}, {12'sd1726, 11'sd716, 13'sd-2231}, {11'sd853, 12'sd-1912, 12'sd1798}},
{{11'sd-834, 11'sd-801, 12'sd1390}, {10'sd420, 11'sd-573, 11'sd-857}, {10'sd-487, 12'sd-1182, 11'sd715}},
{{11'sd-822, 12'sd1732, 10'sd-351}, {11'sd-705, 13'sd2058, 10'sd-420}, {12'sd1917, 12'sd-1293, 12'sd1119}},
{{10'sd276, 9'sd-228, 13'sd2360}, {13'sd-2354, 12'sd1375, 9'sd-222}, {13'sd-3236, 12'sd-1050, 13'sd-2099}},
{{13'sd2094, 12'sd1591, 13'sd-3511}, {12'sd1373, 13'sd2072, 11'sd979}, {11'sd-741, 11'sd-798, 11'sd617}}},
{
{{13'sd2140, 9'sd203, 13'sd2706}, {12'sd1094, 12'sd1739, 10'sd-353}, {12'sd1551, 13'sd-2964, 12'sd1989}},
{{12'sd1732, 13'sd2129, 12'sd1094}, {9'sd154, 13'sd2174, 13'sd2432}, {11'sd869, 5'sd9, 12'sd1148}},
{{13'sd2399, 10'sd-414, 12'sd1635}, {13'sd-2623, 11'sd-914, 12'sd-1326}, {12'sd1312, 12'sd1351, 12'sd-1082}},
{{12'sd1134, 11'sd867, 9'sd-134}, {13'sd-2096, 13'sd-2643, 13'sd2276}, {12'sd1180, 8'sd104, 10'sd428}},
{{11'sd622, 8'sd107, 11'sd844}, {12'sd1154, 10'sd266, 13'sd2243}, {12'sd-1852, 12'sd1189, 12'sd1713}},
{{12'sd1131, 12'sd1879, 12'sd-1339}, {12'sd1405, 13'sd-2279, 12'sd-1769}, {9'sd206, 12'sd1948, 9'sd170}},
{{11'sd782, 12'sd-1076, 13'sd-2144}, {11'sd668, 13'sd2595, 12'sd-1172}, {12'sd1322, 13'sd2140, 13'sd2931}},
{{10'sd274, 11'sd-588, 10'sd297}, {13'sd-2357, 13'sd2246, 12'sd1365}, {12'sd1397, 12'sd1670, 12'sd-1309}},
{{12'sd1428, 13'sd-2464, 12'sd-2023}, {13'sd-2344, 13'sd2291, 11'sd574}, {11'sd-861, 12'sd1117, 11'sd-849}},
{{12'sd1185, 11'sd857, 11'sd-742}, {12'sd-1732, 9'sd-190, 12'sd-1878}, {12'sd1114, 12'sd-1081, 13'sd-2070}},
{{10'sd399, 13'sd-3090, 13'sd2856}, {9'sd-183, 12'sd-1887, 13'sd2121}, {12'sd-1376, 12'sd1932, 13'sd2334}},
{{9'sd-223, 12'sd1554, 13'sd2151}, {13'sd2566, 13'sd2769, 10'sd-325}, {12'sd-1770, 13'sd-2534, 12'sd1295}},
{{11'sd935, 9'sd250, 13'sd-2739}, {12'sd-1906, 13'sd2790, 12'sd1500}, {13'sd3864, 10'sd-417, 11'sd917}},
{{7'sd40, 12'sd-1646, 13'sd2083}, {3'sd-2, 12'sd-1328, 10'sd-481}, {13'sd2402, 13'sd2419, 10'sd288}},
{{13'sd-2122, 12'sd1424, 10'sd477}, {12'sd-1427, 10'sd-474, 12'sd-1618}, {12'sd-2028, 12'sd-1933, 9'sd-138}},
{{13'sd2363, 12'sd1798, 12'sd1030}, {12'sd-1426, 9'sd154, 13'sd3183}, {13'sd2696, 11'sd-615, 12'sd-1885}},
{{12'sd1812, 11'sd601, 11'sd753}, {9'sd-159, 12'sd1463, 13'sd-2140}, {11'sd748, 11'sd-955, 12'sd1068}},
{{12'sd1912, 13'sd2536, 11'sd-826}, {12'sd-1044, 11'sd618, 13'sd-3984}, {11'sd824, 12'sd-1736, 12'sd-1508}},
{{12'sd-1483, 12'sd1240, 12'sd-1140}, {13'sd2143, 13'sd2057, 11'sd627}, {12'sd-1277, 12'sd-1665, 12'sd-1540}},
{{13'sd2086, 13'sd-2614, 10'sd-283}, {12'sd-1926, 12'sd2023, 12'sd1119}, {12'sd-2041, 13'sd2313, 13'sd-2493}},
{{10'sd-395, 13'sd2577, 12'sd1067}, {11'sd1006, 9'sd-130, 11'sd-1015}, {10'sd-473, 12'sd1523, 12'sd-2023}},
{{12'sd-1740, 12'sd-1679, 12'sd-1261}, {13'sd2672, 12'sd1848, 12'sd-1468}, {14'sd4540, 10'sd-477, 13'sd3742}},
{{12'sd1455, 11'sd-863, 12'sd-1190}, {12'sd1607, 12'sd1148, 11'sd615}, {9'sd230, 12'sd1672, 8'sd110}},
{{12'sd1205, 12'sd2038, 11'sd-526}, {11'sd-726, 13'sd-2853, 12'sd1539}, {11'sd1005, 11'sd-568, 11'sd563}},
{{12'sd2007, 13'sd2500, 12'sd-1716}, {11'sd-1006, 13'sd3978, 6'sd19}, {11'sd740, 11'sd-566, 13'sd-2256}},
{{12'sd1032, 8'sd-85, 12'sd1083}, {2'sd-1, 12'sd-1458, 13'sd2733}, {12'sd-2004, 12'sd1414, 12'sd-1049}},
{{12'sd1337, 13'sd2086, 9'sd-207}, {11'sd572, 11'sd-821, 13'sd2419}, {9'sd-154, 12'sd-1527, 12'sd1343}},
{{13'sd-2801, 12'sd1447, 12'sd1127}, {12'sd-1462, 12'sd1244, 13'sd2394}, {12'sd-1707, 4'sd-6, 13'sd2089}},
{{13'sd-3142, 10'sd-425, 11'sd941}, {12'sd-1750, 12'sd-1281, 12'sd-1362}, {7'sd59, 13'sd2094, 11'sd-768}},
{{12'sd1654, 13'sd-2197, 11'sd616}, {12'sd1897, 8'sd-103, 13'sd3200}, {11'sd-884, 12'sd1211, 11'sd572}},
{{13'sd-2563, 11'sd854, 12'sd1846}, {10'sd298, 13'sd-2238, 13'sd-2906}, {11'sd823, 10'sd-261, 13'sd2641}},
{{10'sd340, 10'sd476, 11'sd823}, {12'sd-1057, 13'sd2534, 11'sd705}, {10'sd510, 12'sd-1481, 10'sd401}},
{{13'sd-2358, 12'sd1095, 12'sd1175}, {9'sd-210, 12'sd1600, 11'sd999}, {13'sd-2592, 12'sd1647, 7'sd62}},
{{12'sd1521, 12'sd-1221, 11'sd871}, {10'sd-364, 10'sd501, 13'sd-2126}, {12'sd-1872, 12'sd-1454, 13'sd-2658}},
{{10'sd-346, 11'sd-569, 11'sd1020}, {9'sd161, 12'sd1308, 12'sd1598}, {4'sd-6, 8'sd-75, 13'sd2129}},
{{10'sd-376, 11'sd-911, 12'sd-1903}, {11'sd-946, 10'sd348, 11'sd-534}, {13'sd2529, 12'sd1103, 11'sd732}},
{{9'sd-147, 12'sd1899, 10'sd-445}, {11'sd987, 12'sd1736, 12'sd1914}, {10'sd401, 11'sd1019, 10'sd-311}},
{{10'sd426, 13'sd-2433, 11'sd-837}, {11'sd648, 8'sd-74, 14'sd4234}, {13'sd2901, 12'sd1694, 12'sd1120}},
{{12'sd1816, 11'sd593, 12'sd-1882}, {13'sd3042, 6'sd-16, 7'sd-63}, {12'sd-1105, 9'sd170, 12'sd1825}},
{{12'sd-1045, 9'sd-201, 10'sd388}, {13'sd2668, 9'sd134, 12'sd-1813}, {8'sd78, 11'sd948, 11'sd994}},
{{11'sd530, 13'sd2410, 12'sd1999}, {13'sd2159, 13'sd3152, 9'sd210}, {12'sd1882, 11'sd-874, 12'sd-1998}},
{{13'sd-2055, 11'sd692, 12'sd1784}, {7'sd36, 12'sd-1162, 12'sd-2041}, {13'sd2441, 11'sd-986, 12'sd1321}},
{{11'sd-851, 12'sd-1705, 11'sd693}, {11'sd-787, 12'sd-1359, 12'sd1853}, {11'sd-676, 13'sd2271, 12'sd-1308}},
{{12'sd1682, 11'sd-567, 13'sd2438}, {10'sd-338, 13'sd-2505, 8'sd81}, {12'sd1699, 13'sd-2087, 12'sd1124}},
{{11'sd767, 13'sd-2621, 11'sd608}, {7'sd63, 13'sd-2246, 11'sd-914}, {11'sd-787, 12'sd-1318, 12'sd1322}},
{{11'sd-800, 13'sd-2842, 10'sd-477}, {9'sd254, 10'sd282, 12'sd1654}, {12'sd1648, 12'sd-1543, 10'sd474}},
{{12'sd1378, 12'sd1590, 10'sd323}, {12'sd1664, 8'sd124, 11'sd-941}, {12'sd1091, 12'sd1650, 13'sd2070}},
{{13'sd-2487, 13'sd-2345, 13'sd-2592}, {12'sd-1338, 9'sd161, 11'sd-876}, {11'sd567, 12'sd-1357, 10'sd489}},
{{10'sd362, 9'sd-215, 13'sd2490}, {12'sd1356, 12'sd1287, 13'sd2148}, {12'sd-1632, 11'sd-949, 11'sd-881}},
{{13'sd-2748, 13'sd2535, 12'sd-1863}, {12'sd-1733, 13'sd2204, 13'sd-2222}, {11'sd-912, 12'sd1907, 11'sd-618}},
{{13'sd2075, 11'sd901, 12'sd1212}, {13'sd-2186, 7'sd-33, 11'sd-761}, {13'sd2739, 12'sd1669, 11'sd621}},
{{10'sd481, 12'sd-1656, 13'sd-2480}, {9'sd-150, 12'sd1635, 11'sd-1011}, {12'sd-1618, 9'sd224, 10'sd296}},
{{14'sd4161, 12'sd-1253, 10'sd-365}, {12'sd1123, 10'sd-484, 12'sd1386}, {12'sd-1318, 12'sd1661, 12'sd1457}},
{{12'sd1398, 13'sd-2179, 13'sd-2363}, {11'sd-921, 11'sd833, 13'sd2673}, {10'sd502, 11'sd-909, 4'sd7}},
{{11'sd838, 13'sd2748, 13'sd2402}, {11'sd-801, 10'sd-359, 12'sd1944}, {13'sd2388, 12'sd-1079, 13'sd2903}},
{{11'sd583, 12'sd1704, 9'sd234}, {12'sd-1519, 13'sd-2754, 11'sd-990}, {11'sd-939, 11'sd1001, 12'sd1308}},
{{12'sd1380, 12'sd-1094, 12'sd-1329}, {6'sd-29, 11'sd723, 12'sd1334}, {12'sd2031, 11'sd-726, 12'sd1649}},
{{13'sd3000, 11'sd739, 12'sd-1708}, {13'sd2078, 11'sd623, 9'sd215}, {13'sd-3968, 13'sd-3002, 11'sd-835}},
{{12'sd1526, 13'sd2140, 12'sd1839}, {12'sd-1899, 11'sd-584, 12'sd1229}, {11'sd-694, 12'sd-1831, 10'sd-276}},
{{11'sd-886, 13'sd2694, 12'sd-1488}, {13'sd2273, 9'sd-240, 12'sd1050}, {13'sd2842, 12'sd-1871, 12'sd-1247}},
{{11'sd-625, 11'sd-513, 12'sd-1727}, {12'sd1501, 11'sd-838, 13'sd2605}, {13'sd2292, 13'sd-2965, 10'sd489}},
{{10'sd-475, 11'sd781, 12'sd-1606}, {12'sd1061, 9'sd-169, 13'sd-2299}, {11'sd854, 12'sd-1471, 11'sd572}},
{{12'sd-1034, 12'sd-1564, 10'sd292}, {10'sd-332, 8'sd121, 12'sd1488}, {12'sd1420, 13'sd-2474, 8'sd-102}},
{{10'sd465, 11'sd607, 13'sd3004}, {12'sd-1155, 12'sd1948, 12'sd1691}, {12'sd1763, 13'sd2525, 13'sd2482}}},
{
{{13'sd-2138, 12'sd-1087, 13'sd3268}, {12'sd-1956, 11'sd-763, 12'sd1503}, {13'sd-2153, 12'sd1981, 12'sd1384}},
{{11'sd-700, 13'sd2545, 12'sd-1749}, {12'sd1324, 13'sd2254, 12'sd-1861}, {10'sd-424, 12'sd1664, 9'sd230}},
{{13'sd3168, 12'sd1955, 11'sd-992}, {13'sd2293, 13'sd-2754, 12'sd1691}, {12'sd-1332, 12'sd-1693, 13'sd-3300}},
{{9'sd-167, 9'sd-234, 12'sd-1997}, {12'sd1762, 13'sd-2243, 12'sd1316}, {12'sd1943, 12'sd1231, 12'sd-1989}},
{{12'sd-1684, 12'sd1182, 12'sd-1630}, {12'sd-1113, 9'sd195, 8'sd87}, {12'sd-1767, 13'sd-2957, 12'sd-1532}},
{{10'sd302, 11'sd721, 12'sd-1248}, {12'sd1767, 12'sd1160, 12'sd1113}, {13'sd2702, 12'sd-1283, 13'sd2283}},
{{11'sd-742, 9'sd146, 11'sd823}, {12'sd1347, 10'sd450, 11'sd881}, {11'sd-628, 11'sd582, 12'sd-2043}},
{{9'sd-195, 12'sd2043, 12'sd1179}, {10'sd-497, 11'sd904, 8'sd-90}, {10'sd475, 12'sd-1760, 12'sd1871}},
{{12'sd1889, 12'sd-1977, 9'sd-241}, {12'sd-1055, 10'sd-338, 9'sd-192}, {13'sd2665, 13'sd2355, 12'sd-1578}},
{{12'sd1559, 12'sd1072, 10'sd-361}, {11'sd969, 12'sd1246, 13'sd2796}, {12'sd1323, 11'sd897, 13'sd-2326}},
{{10'sd-342, 10'sd452, 10'sd-415}, {10'sd458, 12'sd-1298, 12'sd-1713}, {8'sd106, 13'sd2117, 12'sd-1174}},
{{12'sd-1538, 11'sd-714, 12'sd1025}, {12'sd1088, 13'sd-2125, 12'sd-1893}, {12'sd-1231, 11'sd-627, 12'sd1353}},
{{8'sd104, 13'sd2458, 12'sd-1659}, {13'sd2391, 12'sd-1313, 12'sd1577}, {13'sd-2227, 12'sd-1847, 13'sd2089}},
{{12'sd1273, 12'sd-1313, 10'sd393}, {13'sd-2602, 13'sd-2686, 12'sd-1705}, {13'sd-2153, 13'sd2506, 13'sd-2222}},
{{11'sd617, 13'sd-2481, 12'sd1757}, {12'sd1630, 13'sd-2258, 13'sd2281}, {8'sd68, 11'sd786, 11'sd642}},
{{10'sd264, 10'sd-289, 11'sd677}, {12'sd1204, 12'sd1049, 12'sd1763}, {9'sd-214, 11'sd-834, 12'sd1563}},
{{11'sd-540, 11'sd673, 11'sd549}, {11'sd-914, 13'sd2194, 11'sd-733}, {11'sd-774, 12'sd-1486, 10'sd-263}},
{{12'sd1481, 13'sd3415, 13'sd2189}, {11'sd669, 13'sd-2858, 13'sd-3648}, {13'sd-2244, 12'sd-1361, 13'sd-3549}},
{{12'sd-1185, 12'sd-1692, 8'sd-94}, {12'sd-2010, 12'sd-1134, 10'sd379}, {12'sd-1303, 13'sd-2487, 13'sd-2364}},
{{12'sd-1723, 11'sd825, 10'sd-420}, {9'sd-182, 13'sd2859, 12'sd1551}, {11'sd-807, 9'sd149, 12'sd-1924}},
{{11'sd612, 9'sd249, 9'sd240}, {13'sd2396, 11'sd-691, 12'sd-1878}, {11'sd-650, 13'sd-2261, 12'sd1985}},
{{11'sd-570, 11'sd579, 12'sd-1316}, {13'sd2246, 12'sd1599, 9'sd161}, {11'sd-554, 12'sd-1919, 12'sd1729}},
{{13'sd2631, 12'sd-1442, 11'sd541}, {11'sd715, 12'sd-1957, 10'sd-411}, {13'sd2533, 11'sd-813, 12'sd-1712}},
{{12'sd-1614, 11'sd636, 11'sd973}, {10'sd332, 11'sd772, 13'sd-2253}, {12'sd1178, 11'sd802, 11'sd914}},
{{11'sd982, 13'sd-2176, 12'sd-1094}, {11'sd628, 12'sd1687, 13'sd-2842}, {13'sd-2087, 13'sd-3016, 13'sd-2296}},
{{12'sd-1654, 12'sd1316, 11'sd640}, {12'sd-1160, 12'sd1219, 11'sd-889}, {11'sd-701, 11'sd-923, 11'sd-713}},
{{11'sd-877, 12'sd1115, 13'sd2715}, {10'sd-256, 10'sd402, 9'sd216}, {12'sd-1913, 13'sd2543, 12'sd2047}},
{{12'sd-1473, 6'sd-29, 10'sd331}, {11'sd850, 12'sd1824, 12'sd1530}, {9'sd-254, 12'sd-1512, 12'sd-1542}},
{{11'sd-688, 13'sd2069, 13'sd2765}, {13'sd2657, 13'sd2157, 12'sd1595}, {10'sd-311, 11'sd-875, 13'sd-2351}},
{{12'sd-1424, 12'sd1894, 12'sd-1925}, {13'sd2521, 13'sd-2367, 12'sd1415}, {13'sd2840, 12'sd1373, 12'sd1974}},
{{10'sd378, 10'sd345, 12'sd1246}, {12'sd-1053, 12'sd-1684, 12'sd1979}, {13'sd2371, 11'sd-842, 11'sd-774}},
{{11'sd-550, 9'sd135, 13'sd-2162}, {12'sd-1394, 12'sd-1540, 11'sd-990}, {10'sd327, 12'sd-1702, 13'sd2148}},
{{12'sd1790, 13'sd-2350, 12'sd2005}, {7'sd-40, 10'sd-359, 12'sd-1932}, {11'sd753, 11'sd-739, 10'sd-363}},
{{13'sd2434, 10'sd-323, 11'sd681}, {13'sd2551, 11'sd515, 13'sd2100}, {12'sd-2029, 13'sd-2236, 12'sd1276}},
{{13'sd-2788, 13'sd2172, 12'sd1607}, {10'sd-399, 12'sd-1540, 12'sd-1630}, {10'sd382, 12'sd-1537, 12'sd1434}},
{{13'sd-2462, 12'sd-1633, 9'sd-204}, {12'sd1468, 12'sd1236, 13'sd-2291}, {11'sd-925, 13'sd2737, 11'sd-1015}},
{{11'sd-741, 13'sd2370, 12'sd-1236}, {10'sd393, 11'sd-1018, 11'sd693}, {13'sd-2681, 12'sd-1250, 11'sd688}},
{{13'sd-3033, 11'sd769, 12'sd-1170}, {11'sd875, 12'sd-1571, 12'sd-1161}, {13'sd-2169, 10'sd-283, 13'sd3101}},
{{13'sd2253, 13'sd-2407, 11'sd727}, {13'sd-3067, 12'sd1336, 8'sd100}, {12'sd1955, 11'sd677, 8'sd124}},
{{13'sd-2440, 11'sd-735, 13'sd2657}, {12'sd-1782, 12'sd-1231, 12'sd2005}, {10'sd-320, 12'sd1764, 13'sd2220}},
{{11'sd733, 11'sd1005, 12'sd-1308}, {12'sd1067, 13'sd2289, 11'sd-975}, {12'sd-1958, 12'sd1096, 12'sd-1875}},
{{12'sd1069, 11'sd-618, 12'sd-1335}, {12'sd1753, 11'sd526, 12'sd1895}, {13'sd2108, 10'sd-509, 13'sd2564}},
{{12'sd1307, 8'sd-120, 12'sd-1106}, {11'sd532, 12'sd-1484, 12'sd1662}, {11'sd956, 9'sd-250, 12'sd-2011}},
{{12'sd-1866, 13'sd-2542, 11'sd-625}, {13'sd-2352, 10'sd-456, 7'sd51}, {12'sd-1758, 10'sd398, 12'sd1451}},
{{13'sd2729, 13'sd-2637, 11'sd584}, {13'sd2595, 8'sd92, 12'sd-1499}, {12'sd1639, 12'sd-1878, 12'sd-1679}},
{{12'sd1448, 13'sd2149, 12'sd1221}, {12'sd1198, 12'sd-1054, 9'sd-142}, {12'sd1884, 12'sd2033, 11'sd753}},
{{11'sd-742, 12'sd1053, 13'sd3240}, {12'sd1549, 13'sd2382, 13'sd2971}, {12'sd-1338, 13'sd-2879, 11'sd-652}},
{{13'sd-2116, 12'sd1183, 10'sd-438}, {13'sd2160, 13'sd-2266, 12'sd-1427}, {13'sd2195, 12'sd-1278, 13'sd-2651}},
{{11'sd-896, 11'sd-839, 12'sd-1270}, {12'sd-1221, 11'sd-577, 12'sd1383}, {12'sd1944, 12'sd-1594, 11'sd-706}},
{{13'sd-2391, 12'sd1080, 13'sd-2645}, {10'sd-462, 11'sd-888, 10'sd-383}, {11'sd-661, 13'sd-2596, 12'sd1391}},
{{9'sd171, 13'sd-2172, 13'sd2341}, {12'sd1486, 13'sd2568, 12'sd1398}, {11'sd701, 12'sd1925, 12'sd-1290}},
{{13'sd2241, 13'sd2155, 10'sd378}, {13'sd2256, 11'sd686, 13'sd-2505}, {11'sd948, 12'sd1551, 12'sd-1026}},
{{13'sd3776, 9'sd-140, 13'sd2883}, {12'sd-2040, 9'sd-253, 11'sd689}, {8'sd127, 13'sd-4016, 12'sd1103}},
{{9'sd-128, 9'sd-247, 12'sd-2033}, {11'sd-779, 13'sd2615, 11'sd907}, {11'sd668, 9'sd-205, 12'sd1347}},
{{12'sd-1112, 11'sd-1003, 8'sd88}, {12'sd1091, 12'sd-1655, 12'sd-1299}, {12'sd1271, 13'sd2649, 12'sd1974}},
{{12'sd1852, 12'sd1124, 10'sd-362}, {12'sd1369, 13'sd2946, 13'sd2638}, {12'sd1616, 11'sd-778, 10'sd-333}},
{{12'sd1240, 13'sd-2067, 12'sd1266}, {8'sd-118, 13'sd2577, 12'sd1319}, {6'sd19, 13'sd-2621, 13'sd-3117}},
{{12'sd1878, 12'sd1163, 13'sd2886}, {12'sd1330, 9'sd-165, 12'sd2028}, {11'sd654, 11'sd-1001, 7'sd-44}},
{{12'sd-1322, 13'sd2264, 12'sd-1129}, {12'sd-1812, 12'sd-1960, 12'sd1866}, {13'sd-2563, 12'sd1884, 12'sd-1726}},
{{11'sd-733, 13'sd2691, 10'sd342}, {12'sd1516, 11'sd-634, 13'sd-2376}, {11'sd-539, 12'sd-1135, 12'sd1875}},
{{12'sd-1171, 13'sd-2289, 12'sd-2038}, {13'sd-2205, 13'sd2176, 13'sd-2503}, {10'sd416, 12'sd-1452, 9'sd158}},
{{10'sd486, 11'sd-807, 12'sd1561}, {13'sd2745, 13'sd2651, 4'sd-7}, {11'sd-804, 13'sd2773, 11'sd-542}},
{{11'sd1022, 7'sd50, 11'sd-781}, {12'sd2046, 12'sd1538, 13'sd-2320}, {12'sd-1026, 12'sd-1662, 11'sd-834}},
{{12'sd1428, 13'sd3190, 12'sd-1317}, {10'sd300, 13'sd2519, 11'sd943}, {12'sd-1173, 9'sd250, 12'sd1509}}},
{
{{13'sd-2686, 11'sd903, 11'sd-643}, {8'sd77, 12'sd-1242, 13'sd2350}, {13'sd-3474, 12'sd-1325, 13'sd2288}},
{{8'sd70, 13'sd2342, 12'sd1712}, {10'sd380, 13'sd3114, 10'sd333}, {10'sd-454, 11'sd-661, 12'sd1509}},
{{3'sd-2, 13'sd2483, 13'sd-2159}, {10'sd-454, 11'sd-804, 11'sd-975}, {13'sd-3742, 12'sd-1156, 14'sd-4118}},
{{13'sd-2475, 12'sd1547, 8'sd103}, {11'sd-601, 13'sd-2110, 12'sd1412}, {13'sd2417, 12'sd1248, 12'sd1390}},
{{13'sd2859, 13'sd2215, 13'sd3286}, {12'sd1085, 12'sd1931, 11'sd-517}, {12'sd1410, 9'sd-184, 12'sd-2011}},
{{13'sd-2139, 12'sd-1911, 11'sd-643}, {12'sd-1558, 13'sd2317, 9'sd-173}, {13'sd-2666, 8'sd-115, 12'sd-1932}},
{{11'sd839, 12'sd-1220, 12'sd1994}, {13'sd-2321, 8'sd-80, 11'sd-825}, {13'sd3050, 9'sd202, 12'sd-1586}},
{{8'sd-85, 11'sd-529, 12'sd-1095}, {12'sd1791, 11'sd-658, 13'sd-2725}, {10'sd-295, 8'sd-90, 13'sd2255}},
{{13'sd-2113, 12'sd1603, 10'sd-511}, {12'sd2030, 13'sd-2349, 12'sd1484}, {13'sd-2494, 13'sd-2905, 10'sd-340}},
{{12'sd2012, 10'sd435, 11'sd861}, {12'sd-1475, 11'sd-889, 12'sd-1570}, {13'sd-2079, 11'sd-978, 11'sd-740}},
{{12'sd1179, 12'sd1989, 13'sd2545}, {12'sd1680, 13'sd2309, 12'sd1976}, {12'sd1285, 14'sd4581, 12'sd1279}},
{{11'sd762, 12'sd1731, 13'sd-2405}, {8'sd-123, 12'sd1844, 13'sd2164}, {13'sd2068, 13'sd-2048, 10'sd-472}},
{{11'sd-968, 13'sd2675, 13'sd-3468}, {13'sd3863, 12'sd-1697, 13'sd-3964}, {12'sd1443, 13'sd3824, 12'sd1174}},
{{13'sd-2285, 8'sd-81, 11'sd-836}, {9'sd197, 12'sd1711, 9'sd-213}, {11'sd-712, 13'sd2629, 12'sd1873}},
{{12'sd1229, 12'sd1324, 12'sd2009}, {12'sd-2042, 13'sd-2075, 12'sd-1829}, {11'sd-622, 8'sd105, 11'sd-967}},
{{11'sd-974, 13'sd2412, 11'sd-923}, {13'sd3671, 13'sd-2724, 13'sd2213}, {13'sd3818, 7'sd-53, 12'sd1206}},
{{11'sd-607, 12'sd1851, 7'sd42}, {12'sd1411, 10'sd-427, 9'sd226}, {13'sd2299, 12'sd1048, 13'sd2796}},
{{12'sd1243, 10'sd-259, 11'sd752}, {12'sd-1858, 11'sd-884, 12'sd-1251}, {14'sd-6146, 11'sd-751, 12'sd-1165}},
{{11'sd974, 12'sd1358, 12'sd1665}, {8'sd105, 10'sd-511, 13'sd-2656}, {13'sd2260, 12'sd-1258, 11'sd-537}},
{{13'sd2180, 12'sd1411, 12'sd1280}, {12'sd1840, 9'sd129, 10'sd388}, {12'sd1100, 11'sd767, 13'sd2322}},
{{11'sd-1013, 13'sd-2603, 13'sd-2150}, {12'sd-1774, 13'sd2713, 12'sd-1931}, {12'sd-1823, 11'sd564, 12'sd-1458}},
{{10'sd423, 8'sd-76, 11'sd968}, {13'sd2941, 12'sd-1151, 12'sd1760}, {13'sd3870, 13'sd-2091, 12'sd-1795}},
{{12'sd-1145, 13'sd2242, 11'sd-814}, {10'sd386, 13'sd2063, 11'sd-858}, {10'sd-301, 13'sd2256, 12'sd1539}},
{{11'sd-817, 13'sd-2080, 12'sd-1902}, {11'sd-529, 12'sd-1740, 12'sd1760}, {11'sd-605, 10'sd275, 12'sd-1045}},
{{11'sd-628, 12'sd-1324, 8'sd86}, {12'sd-1190, 12'sd1428, 12'sd-1237}, {13'sd-2600, 11'sd-812, 13'sd-2217}},
{{12'sd-1676, 9'sd-218, 13'sd2289}, {13'sd2111, 11'sd726, 12'sd-1585}, {12'sd1432, 12'sd1619, 12'sd-1071}},
{{11'sd1017, 11'sd1022, 11'sd750}, {12'sd-1731, 10'sd-470, 12'sd1728}, {13'sd-2804, 12'sd-1954, 13'sd-2675}},
{{11'sd-598, 13'sd2480, 11'sd-529}, {10'sd473, 9'sd-221, 9'sd-217}, {13'sd2413, 12'sd1286, 11'sd-887}},
{{5'sd-11, 13'sd2458, 13'sd2367}, {12'sd1526, 11'sd-814, 12'sd-1299}, {11'sd611, 12'sd-1930, 12'sd-1122}},
{{12'sd-1457, 8'sd93, 12'sd-1721}, {13'sd2986, 13'sd2605, 13'sd2540}, {13'sd3874, 12'sd1563, 12'sd1736}},
{{11'sd-891, 12'sd-1707, 11'sd-554}, {12'sd1498, 12'sd1091, 13'sd2980}, {8'sd125, 13'sd2279, 13'sd-2232}},
{{12'sd-1192, 13'sd3135, 12'sd2042}, {13'sd-2472, 13'sd-2511, 11'sd-631}, {11'sd-938, 11'sd-533, 12'sd-2029}},
{{8'sd-70, 13'sd-2148, 12'sd-1560}, {10'sd474, 12'sd-1567, 12'sd-1589}, {12'sd-1100, 11'sd-550, 13'sd-2294}},
{{12'sd-1371, 13'sd2499, 13'sd-2274}, {11'sd-672, 12'sd1909, 13'sd2117}, {11'sd620, 13'sd2538, 12'sd-1478}},
{{13'sd-3209, 13'sd-2503, 12'sd1874}, {12'sd-1196, 10'sd-327, 5'sd-13}, {10'sd-462, 9'sd163, 13'sd2913}},
{{12'sd-1362, 12'sd-1751, 13'sd-2567}, {12'sd1995, 12'sd1700, 12'sd1706}, {11'sd-525, 12'sd1185, 12'sd1451}},
{{13'sd-2536, 12'sd1775, 12'sd-1360}, {12'sd1567, 12'sd1502, 11'sd-981}, {13'sd-2538, 12'sd-1323, 10'sd-431}},
{{10'sd362, 12'sd2006, 11'sd918}, {14'sd4389, 12'sd-1721, 13'sd2301}, {10'sd506, 14'sd-4135, 9'sd179}},
{{11'sd-808, 13'sd2258, 13'sd2627}, {11'sd574, 10'sd-278, 12'sd1339}, {13'sd2973, 12'sd2043, 12'sd-1304}},
{{12'sd1506, 11'sd722, 11'sd792}, {13'sd2871, 10'sd-444, 11'sd-552}, {13'sd-2392, 13'sd-2902, 10'sd284}},
{{13'sd2112, 13'sd2736, 8'sd-89}, {11'sd-669, 13'sd2310, 11'sd-728}, {12'sd1051, 11'sd517, 13'sd-2698}},
{{9'sd-229, 12'sd-1462, 12'sd1729}, {11'sd580, 13'sd-2551, 12'sd1765}, {12'sd-1990, 11'sd640, 12'sd-1355}},
{{11'sd801, 11'sd-784, 12'sd1544}, {13'sd-2310, 10'sd-413, 12'sd-1810}, {12'sd-1898, 13'sd2588, 13'sd3190}},
{{13'sd-2639, 13'sd2190, 13'sd-2884}, {13'sd-2241, 10'sd-474, 11'sd-701}, {8'sd98, 14'sd4499, 13'sd2213}},
{{13'sd-2527, 13'sd2229, 11'sd-868}, {12'sd-1836, 11'sd619, 12'sd-1729}, {12'sd1650, 13'sd2111, 12'sd-1110}},
{{9'sd231, 12'sd-1226, 12'sd-1705}, {13'sd-2852, 11'sd726, 12'sd1853}, {8'sd-71, 13'sd-2801, 11'sd821}},
{{10'sd384, 12'sd1257, 12'sd1840}, {11'sd-657, 10'sd-374, 10'sd301}, {9'sd-197, 12'sd-1187, 13'sd2608}},
{{11'sd-744, 10'sd-368, 12'sd-1700}, {13'sd2068, 12'sd-1083, 12'sd-1822}, {11'sd-811, 12'sd-1537, 10'sd423}},
{{10'sd349, 11'sd973, 13'sd-2137}, {13'sd-2406, 13'sd-2438, 12'sd-1675}, {12'sd-1266, 12'sd-1037, 12'sd1682}},
{{12'sd1366, 12'sd-1140, 13'sd2305}, {11'sd691, 12'sd-1393, 12'sd1472}, {13'sd-2211, 10'sd311, 9'sd139}},
{{6'sd-24, 9'sd131, 12'sd-1401}, {11'sd686, 12'sd-1207, 12'sd1933}, {13'sd2988, 11'sd-809, 13'sd-2342}},
{{12'sd-1829, 12'sd-1622, 12'sd1309}, {12'sd-1293, 12'sd1921, 11'sd901}, {10'sd-484, 11'sd-539, 11'sd835}},
{{11'sd-561, 11'sd1016, 14'sd4696}, {12'sd-1881, 9'sd-210, 11'sd581}, {12'sd-2013, 13'sd-3249, 11'sd-712}},
{{11'sd-942, 11'sd863, 13'sd-2295}, {6'sd21, 10'sd508, 10'sd472}, {12'sd-1246, 13'sd-2207, 12'sd-1968}},
{{12'sd-1678, 13'sd2088, 12'sd-1251}, {12'sd1490, 10'sd389, 10'sd-493}, {9'sd-137, 12'sd1528, 12'sd-1954}},
{{11'sd771, 12'sd1941, 13'sd2127}, {12'sd2028, 12'sd-1078, 12'sd1982}, {13'sd-3068, 10'sd335, 11'sd1017}},
{{13'sd-3113, 11'sd675, 12'sd-1272}, {13'sd2661, 11'sd-874, 10'sd-339}, {11'sd555, 10'sd-494, 12'sd1717}},
{{13'sd3027, 14'sd4611, 13'sd3515}, {13'sd-3396, 9'sd-249, 13'sd-3962}, {14'sd-5285, 13'sd-3819, 12'sd-2029}},
{{11'sd-944, 9'sd-131, 13'sd-2103}, {11'sd868, 10'sd-457, 13'sd-3694}, {11'sd-857, 13'sd2439, 7'sd-43}},
{{12'sd-1846, 12'sd-1689, 12'sd-1777}, {13'sd2566, 12'sd-1758, 11'sd-831}, {12'sd1720, 10'sd317, 10'sd323}},
{{13'sd2862, 12'sd-1687, 12'sd-1428}, {11'sd-602, 12'sd-1837, 13'sd-3071}, {13'sd2896, 13'sd-2439, 12'sd1840}},
{{12'sd1550, 13'sd-2381, 12'sd-1930}, {12'sd-1848, 9'sd-219, 12'sd-1509}, {13'sd2412, 11'sd821, 13'sd2301}},
{{12'sd-1810, 11'sd736, 13'sd-2837}, {13'sd-2481, 12'sd1121, 13'sd3064}, {13'sd-2202, 12'sd1418, 10'sd311}},
{{13'sd2074, 12'sd-1267, 11'sd-629}, {12'sd1480, 10'sd-307, 12'sd-1949}, {13'sd-2750, 13'sd-3566, 13'sd-2306}}},
{
{{13'sd-2745, 13'sd-3049, 13'sd-3731}, {11'sd890, 11'sd548, 14'sd-4231}, {12'sd1540, 13'sd2703, 12'sd1352}},
{{13'sd-2127, 11'sd719, 13'sd-2692}, {13'sd-2607, 11'sd665, 9'sd152}, {12'sd-1532, 6'sd-17, 11'sd682}},
{{9'sd135, 9'sd-211, 13'sd-2898}, {12'sd-1154, 13'sd-2224, 13'sd-2992}, {12'sd-1909, 10'sd-318, 10'sd344}},
{{13'sd2481, 13'sd-2646, 12'sd1492}, {13'sd2578, 13'sd2236, 13'sd2445}, {12'sd1823, 12'sd-1841, 11'sd649}},
{{13'sd2835, 13'sd-2930, 12'sd-1775}, {12'sd1479, 12'sd-1714, 13'sd2125}, {12'sd-1101, 12'sd-1410, 12'sd1530}},
{{12'sd2031, 13'sd-2137, 12'sd1530}, {11'sd-741, 12'sd1925, 12'sd-1575}, {12'sd1258, 11'sd1015, 13'sd2815}},
{{10'sd266, 12'sd1920, 13'sd-2507}, {11'sd836, 8'sd-98, 12'sd1237}, {13'sd-2654, 10'sd-355, 11'sd-737}},
{{11'sd-644, 13'sd-2410, 12'sd-1875}, {12'sd-1497, 13'sd-2116, 11'sd558}, {13'sd2145, 9'sd167, 9'sd-196}},
{{10'sd430, 13'sd-2452, 9'sd250}, {12'sd1818, 12'sd1480, 13'sd2470}, {12'sd2043, 12'sd-1187, 13'sd-2659}},
{{13'sd-2384, 12'sd-2042, 13'sd3016}, {13'sd-2790, 12'sd-1258, 7'sd62}, {12'sd1390, 12'sd1253, 10'sd-502}},
{{10'sd-478, 13'sd2553, 13'sd2848}, {13'sd-2679, 12'sd1398, 12'sd1551}, {13'sd-3120, 12'sd1035, 10'sd510}},
{{12'sd-1844, 10'sd-295, 6'sd-30}, {11'sd854, 11'sd651, 12'sd-1671}, {10'sd-452, 12'sd-1875, 10'sd-500}},
{{11'sd-677, 13'sd2122, 13'sd-2333}, {12'sd2045, 10'sd-292, 11'sd540}, {11'sd-866, 13'sd-2816, 12'sd-1302}},
{{13'sd2548, 11'sd550, 12'sd1254}, {12'sd-1576, 13'sd-2712, 13'sd-2540}, {11'sd-793, 10'sd-412, 13'sd2630}},
{{11'sd687, 10'sd-423, 13'sd2493}, {11'sd-560, 11'sd792, 12'sd1132}, {12'sd-1970, 12'sd-1629, 12'sd1271}},
{{12'sd-1330, 10'sd-271, 11'sd889}, {12'sd1367, 12'sd-1877, 11'sd595}, {10'sd-334, 10'sd429, 9'sd234}},
{{7'sd-45, 12'sd-1877, 12'sd1903}, {13'sd3229, 12'sd-1430, 12'sd1487}, {13'sd2185, 10'sd-399, 12'sd-1471}},
{{11'sd-984, 13'sd2815, 14'sd4389}, {12'sd-1965, 7'sd62, 13'sd3826}, {13'sd-2334, 13'sd2939, 12'sd1298}},
{{10'sd286, 12'sd-1172, 13'sd-2281}, {12'sd1061, 11'sd918, 10'sd-301}, {8'sd76, 11'sd540, 13'sd2626}},
{{13'sd-2603, 10'sd-393, 11'sd728}, {12'sd1117, 12'sd-1969, 11'sd-826}, {9'sd238, 11'sd538, 10'sd-259}},
{{12'sd-1577, 11'sd712, 12'sd-1103}, {13'sd2385, 12'sd-1360, 7'sd-50}, {12'sd-1871, 13'sd-2769, 12'sd1231}},
{{12'sd-1937, 12'sd-1406, 13'sd-3106}, {12'sd1643, 11'sd695, 10'sd387}, {13'sd-2733, 11'sd535, 13'sd-2520}},
{{4'sd6, 12'sd1551, 12'sd1127}, {13'sd-2511, 11'sd-588, 6'sd-21}, {12'sd-1688, 12'sd-1087, 12'sd-1997}},
{{10'sd354, 13'sd2654, 10'sd-381}, {13'sd-2519, 8'sd103, 12'sd1330}, {11'sd687, 13'sd-2565, 13'sd-2937}},
{{13'sd-2612, 10'sd379, 13'sd-3158}, {10'sd348, 12'sd-1459, 11'sd583}, {10'sd324, 12'sd1560, 12'sd-1313}},
{{13'sd2772, 11'sd977, 12'sd-1597}, {13'sd-2079, 12'sd-1201, 12'sd1662}, {11'sd-527, 12'sd-1562, 12'sd1374}},
{{10'sd468, 13'sd-2472, 12'sd-1317}, {11'sd595, 12'sd1874, 12'sd-1063}, {11'sd700, 10'sd-401, 12'sd1579}},
{{13'sd2510, 11'sd-1015, 12'sd1493}, {11'sd-891, 12'sd1557, 12'sd2011}, {7'sd-32, 11'sd-666, 12'sd-1853}},
{{13'sd2730, 10'sd-418, 13'sd2696}, {11'sd-996, 11'sd735, 12'sd2037}, {13'sd2079, 10'sd261, 13'sd2693}},
{{12'sd-1939, 11'sd526, 12'sd1777}, {9'sd250, 12'sd1651, 9'sd216}, {9'sd207, 9'sd-161, 13'sd-2086}},
{{12'sd-1657, 11'sd555, 11'sd-745}, {12'sd-1936, 12'sd1745, 11'sd-727}, {13'sd-2140, 12'sd1526, 10'sd278}},
{{12'sd1593, 12'sd1389, 12'sd1037}, {13'sd3429, 13'sd2187, 12'sd1879}, {12'sd1120, 12'sd1339, 13'sd-3507}},
{{13'sd2236, 12'sd-1284, 11'sd-812}, {13'sd-2455, 12'sd1157, 12'sd1783}, {12'sd-1551, 13'sd-2354, 12'sd-1628}},
{{11'sd-583, 8'sd86, 11'sd897}, {12'sd-1971, 13'sd2556, 10'sd466}, {9'sd251, 13'sd-2346, 9'sd230}},
{{12'sd1706, 12'sd1753, 13'sd-3153}, {11'sd645, 9'sd150, 10'sd-351}, {9'sd249, 11'sd-706, 11'sd879}},
{{13'sd2695, 3'sd2, 12'sd-1488}, {11'sd-716, 11'sd-758, 13'sd-2442}, {10'sd-509, 12'sd1516, 10'sd470}},
{{11'sd573, 10'sd-451, 12'sd1114}, {12'sd-1470, 12'sd1113, 12'sd1087}, {13'sd2219, 12'sd-1631, 13'sd-2282}},
{{13'sd2734, 11'sd-986, 8'sd-114}, {10'sd436, 13'sd2429, 9'sd-196}, {13'sd3162, 13'sd2913, 11'sd593}},
{{11'sd720, 10'sd-399, 12'sd-1331}, {12'sd1287, 8'sd127, 11'sd-678}, {10'sd-470, 1'sd0, 13'sd3098}},
{{12'sd1171, 11'sd-515, 11'sd868}, {12'sd1125, 12'sd-1060, 10'sd288}, {10'sd446, 9'sd210, 13'sd2866}},
{{11'sd-988, 11'sd675, 8'sd-110}, {12'sd-1032, 12'sd-1804, 13'sd2391}, {13'sd-2993, 10'sd-405, 12'sd1733}},
{{12'sd-1381, 11'sd-961, 11'sd664}, {10'sd-291, 9'sd167, 9'sd175}, {12'sd2030, 10'sd-369, 9'sd-242}},
{{10'sd-339, 10'sd279, 11'sd-924}, {13'sd-2049, 12'sd-1101, 12'sd1558}, {7'sd-40, 13'sd-2099, 13'sd-2448}},
{{13'sd2750, 13'sd-2642, 13'sd3003}, {11'sd874, 11'sd516, 12'sd1158}, {13'sd2828, 11'sd925, 10'sd-441}},
{{12'sd-1628, 13'sd2508, 8'sd66}, {13'sd-2745, 11'sd871, 9'sd-183}, {13'sd-2234, 11'sd-772, 13'sd2482}},
{{12'sd-1964, 12'sd1061, 12'sd1322}, {12'sd-1339, 10'sd304, 13'sd2221}, {11'sd-520, 13'sd-2194, 8'sd-73}},
{{12'sd1822, 13'sd2900, 13'sd-2452}, {12'sd-1261, 12'sd-1882, 10'sd450}, {12'sd1093, 9'sd-180, 12'sd2036}},
{{12'sd-1619, 12'sd-1505, 12'sd1316}, {10'sd-494, 11'sd-596, 11'sd-835}, {12'sd-1251, 12'sd1866, 12'sd-1381}},
{{13'sd2614, 13'sd-2415, 12'sd1698}, {10'sd-422, 12'sd1783, 11'sd-995}, {11'sd713, 11'sd-871, 11'sd-543}},
{{12'sd-2018, 11'sd-678, 13'sd-2092}, {13'sd-2168, 9'sd-210, 13'sd-2332}, {10'sd-334, 12'sd1933, 10'sd479}},
{{12'sd1165, 13'sd-2066, 10'sd-426}, {12'sd-1299, 12'sd1639, 13'sd-2057}, {11'sd-865, 10'sd-375, 13'sd2788}},
{{13'sd-2191, 9'sd157, 10'sd389}, {9'sd231, 13'sd-2983, 10'sd303}, {12'sd1871, 12'sd-2042, 12'sd1884}},
{{13'sd-2193, 14'sd4316, 13'sd3994}, {12'sd-1337, 13'sd3097, 14'sd4715}, {12'sd1869, 12'sd1670, 10'sd-348}},
{{12'sd-1097, 12'sd1535, 11'sd-812}, {11'sd-966, 12'sd-1394, 12'sd1517}, {11'sd600, 13'sd2955, 13'sd-2235}},
{{8'sd-97, 11'sd1005, 12'sd1871}, {11'sd943, 10'sd-479, 12'sd-1864}, {10'sd405, 12'sd-1252, 10'sd452}},
{{12'sd1808, 11'sd-829, 11'sd707}, {8'sd70, 13'sd2300, 11'sd-969}, {10'sd495, 13'sd-2182, 13'sd-2052}},
{{13'sd-2696, 12'sd-1770, 13'sd2871}, {8'sd-74, 12'sd1209, 12'sd-1050}, {8'sd107, 10'sd-492, 13'sd2558}},
{{12'sd1879, 11'sd-835, 13'sd2778}, {14'sd4156, 12'sd-1188, 12'sd1227}, {12'sd1549, 13'sd2546, 12'sd-1596}},
{{13'sd3775, 12'sd1556, 12'sd1792}, {13'sd2408, 7'sd-48, 12'sd-1205}, {10'sd276, 12'sd-1648, 14'sd-4163}},
{{11'sd699, 12'sd-1822, 10'sd-327}, {11'sd949, 12'sd-1138, 10'sd376}, {13'sd2060, 11'sd-885, 12'sd-1682}},
{{12'sd1751, 13'sd-2886, 12'sd-1104}, {12'sd-1495, 13'sd-2516, 11'sd888}, {11'sd-588, 13'sd-2214, 13'sd-3022}},
{{12'sd1578, 11'sd-572, 13'sd2351}, {13'sd-2174, 12'sd1600, 12'sd-1108}, {12'sd1083, 12'sd-1566, 12'sd-1735}},
{{13'sd2064, 12'sd1859, 11'sd-678}, {10'sd-394, 13'sd2317, 13'sd2347}, {12'sd-1208, 11'sd-623, 12'sd1744}},
{{12'sd-1718, 13'sd-2607, 13'sd-3331}, {12'sd-1430, 13'sd-2328, 13'sd-2875}, {11'sd836, 13'sd2075, 10'sd-440}}},
{
{{12'sd1531, 12'sd1562, 11'sd-633}, {11'sd702, 13'sd-3803, 9'sd-153}, {13'sd2669, 13'sd3891, 13'sd3825}},
{{12'sd1413, 9'sd-246, 10'sd-481}, {13'sd2734, 13'sd2168, 12'sd1892}, {13'sd-2185, 7'sd-57, 11'sd-818}},
{{11'sd-980, 12'sd-1217, 13'sd2936}, {11'sd-702, 8'sd-84, 8'sd-87}, {10'sd505, 12'sd1232, 8'sd-124}},
{{13'sd-2076, 12'sd1180, 10'sd-268}, {12'sd1736, 12'sd-2022, 13'sd-3469}, {12'sd1361, 12'sd-1119, 11'sd-1018}},
{{13'sd3686, 13'sd-3072, 13'sd-2840}, {10'sd-466, 12'sd-1243, 11'sd-589}, {13'sd2613, 6'sd21, 13'sd-2145}},
{{12'sd-2026, 11'sd773, 11'sd978}, {12'sd-1841, 11'sd-537, 12'sd1909}, {11'sd682, 11'sd790, 12'sd-1049}},
{{8'sd-81, 12'sd-1427, 11'sd556}, {9'sd148, 13'sd2804, 13'sd3114}, {13'sd-2919, 11'sd620, 12'sd-1640}},
{{11'sd-834, 12'sd-1259, 11'sd619}, {10'sd-485, 13'sd-3208, 10'sd-511}, {10'sd-352, 13'sd-3556, 12'sd-1729}},
{{13'sd2213, 12'sd1467, 12'sd1515}, {12'sd1442, 13'sd2263, 12'sd-1957}, {8'sd105, 12'sd-1160, 12'sd1425}},
{{13'sd2540, 13'sd-2111, 13'sd-2505}, {12'sd1769, 13'sd-3726, 13'sd2500}, {13'sd2524, 9'sd189, 11'sd-651}},
{{14'sd-4118, 13'sd-2656, 14'sd-4102}, {13'sd-3913, 12'sd1860, 10'sd290}, {12'sd-2007, 13'sd-2543, 11'sd-729}},
{{11'sd-902, 13'sd-2121, 13'sd-2822}, {11'sd-885, 11'sd-700, 13'sd-3036}, {12'sd-1123, 10'sd-453, 11'sd-653}},
{{13'sd-2173, 12'sd1874, 13'sd3796}, {11'sd910, 9'sd-132, 13'sd2684}, {13'sd-4055, 12'sd-1956, 12'sd-1386}},
{{12'sd1466, 10'sd321, 12'sd1658}, {13'sd-2692, 12'sd-1920, 13'sd-2320}, {12'sd1082, 10'sd300, 9'sd221}},
{{11'sd-861, 12'sd1864, 9'sd166}, {13'sd2260, 9'sd141, 12'sd1524}, {12'sd-1566, 12'sd-1525, 12'sd1721}},
{{11'sd-944, 13'sd-2125, 13'sd2588}, {13'sd2243, 9'sd-157, 11'sd-706}, {13'sd2761, 8'sd86, 13'sd-3878}},
{{12'sd-1196, 9'sd199, 12'sd1931}, {8'sd119, 10'sd-258, 13'sd2749}, {13'sd-2395, 13'sd-2189, 13'sd-2224}},
{{14'sd5046, 13'sd2712, 9'sd-198}, {12'sd1760, 14'sd-4257, 12'sd1882}, {10'sd-395, 12'sd-1993, 13'sd-2165}},
{{12'sd1127, 13'sd-2846, 12'sd-1738}, {10'sd298, 12'sd1054, 12'sd1683}, {11'sd634, 11'sd522, 13'sd-3163}},
{{9'sd168, 10'sd-432, 13'sd3259}, {13'sd-2569, 12'sd1400, 13'sd3219}, {13'sd-3802, 14'sd-4262, 13'sd-2250}},
{{12'sd-1112, 10'sd276, 12'sd1381}, {11'sd-649, 12'sd-2036, 12'sd1991}, {12'sd-1509, 12'sd-1976, 10'sd-480}},
{{12'sd1579, 12'sd1051, 11'sd898}, {14'sd4537, 12'sd1723, 13'sd2795}, {13'sd2859, 9'sd206, 12'sd-1626}},
{{13'sd-2612, 7'sd-33, 11'sd536}, {13'sd-2667, 12'sd1858, 11'sd-744}, {11'sd-545, 13'sd2349, 12'sd1535}},
{{10'sd315, 12'sd-2036, 11'sd627}, {12'sd1931, 8'sd-73, 13'sd2552}, {10'sd-363, 9'sd198, 12'sd-1664}},
{{12'sd1442, 9'sd217, 13'sd-2356}, {12'sd1186, 13'sd2244, 12'sd1747}, {13'sd2240, 14'sd4545, 13'sd2154}},
{{13'sd-2994, 10'sd481, 8'sd105}, {13'sd-2739, 6'sd16, 12'sd1447}, {12'sd1250, 12'sd1788, 13'sd-3463}},
{{13'sd2162, 11'sd-769, 11'sd-955}, {12'sd-1309, 10'sd-393, 13'sd-2716}, {11'sd690, 12'sd1440, 12'sd1662}},
{{11'sd951, 12'sd-1253, 10'sd-332}, {12'sd1044, 12'sd-1912, 11'sd-576}, {12'sd-1077, 12'sd1090, 13'sd-3248}},
{{10'sd-387, 14'sd4659, 13'sd2546}, {12'sd-1296, 11'sd-531, 12'sd-1342}, {11'sd-968, 10'sd-501, 12'sd-1905}},
{{12'sd1235, 13'sd2428, 10'sd-467}, {13'sd3777, 13'sd3703, 13'sd3427}, {6'sd-19, 12'sd1530, 13'sd-3279}},
{{12'sd-1533, 13'sd-2429, 13'sd2636}, {13'sd2489, 13'sd2983, 13'sd3230}, {13'sd-3758, 12'sd2037, 12'sd-1804}},
{{13'sd-3275, 13'sd-3690, 12'sd-1413}, {13'sd-3402, 13'sd-3271, 10'sd-268}, {13'sd-2653, 12'sd-1880, 13'sd-3489}},
{{11'sd-821, 13'sd-2269, 9'sd199}, {10'sd-500, 12'sd-1976, 13'sd3526}, {13'sd2098, 11'sd687, 13'sd2129}},
{{13'sd-3012, 11'sd-838, 9'sd-164}, {12'sd1620, 12'sd-1028, 12'sd-1311}, {12'sd-1423, 12'sd-1097, 8'sd97}},
{{6'sd-28, 12'sd1217, 9'sd174}, {13'sd-3616, 12'sd1910, 13'sd-2646}, {10'sd346, 13'sd2403, 10'sd334}},
{{11'sd-599, 13'sd-2112, 11'sd690}, {12'sd-1453, 13'sd2116, 13'sd-3677}, {13'sd2977, 12'sd-2013, 12'sd-1444}},
{{12'sd1982, 13'sd-2080, 13'sd2143}, {12'sd1725, 12'sd-1124, 11'sd522}, {12'sd-1548, 11'sd-661, 13'sd-2381}},
{{8'sd103, 8'sd90, 12'sd1821}, {9'sd153, 11'sd-715, 12'sd-1855}, {13'sd2156, 8'sd82, 13'sd-2243}},
{{13'sd-2263, 12'sd1362, 12'sd1868}, {12'sd1537, 12'sd-1302, 12'sd1069}, {14'sd-5171, 13'sd-2459, 13'sd-3616}},
{{13'sd-3058, 12'sd1576, 14'sd4304}, {13'sd-3502, 12'sd-1439, 12'sd1531}, {12'sd1716, 11'sd-591, 12'sd-1603}},
{{6'sd-27, 12'sd-1223, 9'sd-195}, {12'sd1043, 11'sd-674, 12'sd-1723}, {11'sd755, 12'sd1549, 13'sd-2148}},
{{13'sd3423, 12'sd-1095, 13'sd-2663}, {13'sd2748, 12'sd-1040, 13'sd-2582}, {12'sd1073, 11'sd-540, 12'sd-1553}},
{{12'sd-1212, 12'sd1480, 13'sd-2091}, {12'sd-1026, 13'sd-2156, 10'sd388}, {10'sd-302, 12'sd-1831, 10'sd464}},
{{12'sd-1755, 12'sd1261, 13'sd-2121}, {4'sd-6, 12'sd1423, 12'sd1141}, {12'sd-1268, 10'sd-336, 10'sd382}},
{{8'sd-87, 13'sd3174, 11'sd-551}, {12'sd-1742, 12'sd1893, 12'sd-1030}, {12'sd-1971, 10'sd-432, 9'sd207}},
{{13'sd2401, 11'sd830, 12'sd-1365}, {11'sd-916, 11'sd-839, 12'sd1314}, {12'sd1913, 13'sd2138, 12'sd-1384}},
{{11'sd-614, 11'sd-844, 12'sd1737}, {11'sd-828, 11'sd934, 12'sd-1122}, {12'sd1440, 11'sd-939, 11'sd771}},
{{13'sd2079, 12'sd-1905, 11'sd834}, {8'sd64, 12'sd-1177, 12'sd-1713}, {13'sd2060, 13'sd2471, 11'sd515}},
{{11'sd-688, 12'sd1090, 12'sd-1122}, {12'sd-1897, 13'sd2834, 12'sd-1767}, {11'sd922, 12'sd1925, 12'sd1516}},
{{12'sd-1706, 13'sd2891, 8'sd81}, {13'sd2311, 12'sd1475, 13'sd-2098}, {12'sd-1706, 11'sd629, 11'sd-741}},
{{11'sd-842, 11'sd971, 12'sd-1746}, {11'sd788, 13'sd2488, 13'sd-2631}, {12'sd-1792, 10'sd-500, 13'sd-2474}},
{{12'sd1459, 8'sd-108, 13'sd-2799}, {11'sd937, 12'sd1277, 12'sd-1432}, {12'sd1550, 13'sd2656, 12'sd-1288}},
{{13'sd2323, 9'sd239, 10'sd-449}, {12'sd1889, 13'sd3058, 12'sd1558}, {13'sd3168, 12'sd1865, 12'sd1555}},
{{11'sd649, 12'sd1868, 11'sd858}, {11'sd-976, 6'sd-29, 11'sd621}, {11'sd712, 13'sd-2078, 12'sd-1908}},
{{12'sd-2001, 8'sd-97, 9'sd-171}, {12'sd-1395, 12'sd-1386, 12'sd-1543}, {10'sd-264, 13'sd-2254, 12'sd-1192}},
{{13'sd-2750, 10'sd-295, 10'sd310}, {10'sd426, 13'sd2061, 12'sd1877}, {11'sd532, 12'sd1904, 11'sd-893}},
{{12'sd-1558, 11'sd-692, 11'sd-813}, {12'sd-1072, 10'sd-311, 11'sd836}, {8'sd103, 12'sd-1083, 12'sd1061}},
{{13'sd-3029, 12'sd-1178, 13'sd2903}, {12'sd-1077, 11'sd-611, 13'sd2379}, {10'sd-280, 11'sd-932, 12'sd2013}},
{{6'sd-26, 12'sd-1605, 12'sd1801}, {13'sd-2763, 12'sd-1754, 12'sd-1399}, {13'sd2203, 8'sd126, 12'sd-1607}},
{{9'sd222, 12'sd1389, 7'sd-35}, {12'sd-1219, 10'sd-310, 10'sd-267}, {11'sd-966, 10'sd306, 12'sd-1862}},
{{12'sd-2032, 13'sd-2856, 5'sd-8}, {12'sd-1823, 11'sd997, 12'sd-1199}, {13'sd2804, 13'sd-2432, 12'sd1083}},
{{12'sd1439, 11'sd692, 10'sd-486}, {12'sd1936, 13'sd-2378, 12'sd-1410}, {12'sd1353, 13'sd-2596, 10'sd424}},
{{10'sd-452, 11'sd916, 11'sd-966}, {8'sd-119, 13'sd-2275, 12'sd1371}, {12'sd1389, 12'sd-1160, 12'sd1614}},
{{11'sd659, 13'sd3129, 13'sd2708}, {12'sd1989, 12'sd-1448, 11'sd551}, {13'sd3188, 13'sd3604, 12'sd1525}}},
{
{{13'sd-2198, 12'sd2028, 12'sd-1728}, {13'sd-2467, 11'sd739, 12'sd-1680}, {11'sd-669, 13'sd-2693, 12'sd1780}},
{{13'sd3047, 13'sd-2138, 13'sd-2943}, {10'sd437, 12'sd1450, 12'sd-1743}, {13'sd2142, 4'sd5, 11'sd707}},
{{12'sd-1274, 9'sd175, 10'sd-486}, {12'sd1365, 9'sd-151, 11'sd-538}, {13'sd-2279, 13'sd-2310, 13'sd-3234}},
{{12'sd-2035, 12'sd2026, 13'sd2393}, {13'sd-2753, 13'sd-2779, 13'sd-3012}, {11'sd709, 11'sd855, 12'sd1255}},
{{10'sd355, 13'sd2808, 12'sd-1427}, {12'sd1948, 6'sd-18, 9'sd245}, {13'sd2192, 11'sd-915, 12'sd-1083}},
{{12'sd-1382, 13'sd2763, 13'sd2566}, {13'sd2362, 12'sd1554, 12'sd-1444}, {11'sd793, 12'sd1202, 11'sd512}},
{{12'sd-1962, 13'sd2435, 13'sd-2168}, {10'sd327, 10'sd-291, 12'sd1210}, {11'sd553, 11'sd-866, 12'sd-1515}},
{{9'sd188, 12'sd-1288, 11'sd625}, {13'sd-2078, 13'sd2320, 12'sd1837}, {12'sd-1816, 10'sd277, 13'sd2572}},
{{10'sd-378, 9'sd170, 11'sd-826}, {12'sd1530, 12'sd-2000, 10'sd-357}, {12'sd1064, 11'sd-996, 12'sd1584}},
{{11'sd-873, 12'sd1876, 12'sd-1620}, {13'sd2745, 12'sd-1689, 13'sd-2155}, {10'sd-509, 9'sd-206, 12'sd1555}},
{{14'sd-4595, 13'sd-2922, 9'sd177}, {11'sd-578, 12'sd-1737, 13'sd2794}, {10'sd386, 13'sd2089, 13'sd2557}},
{{12'sd-1683, 10'sd471, 13'sd-2552}, {13'sd-2451, 11'sd-961, 11'sd-1014}, {13'sd2384, 12'sd-1790, 9'sd132}},
{{7'sd-40, 10'sd380, 12'sd-1791}, {11'sd637, 12'sd1217, 12'sd-1406}, {13'sd2496, 12'sd-1298, 13'sd-2068}},
{{13'sd-2420, 11'sd-629, 12'sd1369}, {13'sd-2740, 11'sd536, 12'sd1130}, {11'sd-891, 11'sd-513, 11'sd656}},
{{13'sd-2115, 12'sd-1515, 7'sd-52}, {8'sd-77, 10'sd-457, 13'sd2049}, {12'sd-1619, 12'sd-1734, 13'sd2271}},
{{13'sd-2067, 13'sd-3038, 12'sd1740}, {13'sd2269, 7'sd-61, 13'sd-2770}, {13'sd2578, 11'sd618, 13'sd-2451}},
{{13'sd2644, 11'sd-654, 10'sd-257}, {11'sd613, 11'sd-605, 12'sd-1620}, {12'sd-1217, 12'sd-1703, 10'sd329}},
{{11'sd590, 12'sd1880, 12'sd1969}, {13'sd3352, 13'sd2657, 9'sd173}, {13'sd-3366, 13'sd-3884, 10'sd-268}},
{{11'sd-992, 8'sd-68, 9'sd-171}, {13'sd2166, 10'sd439, 10'sd434}, {12'sd1105, 12'sd-1613, 12'sd1069}},
{{12'sd-1701, 12'sd1996, 10'sd-376}, {12'sd1588, 11'sd632, 13'sd3341}, {12'sd1709, 10'sd377, 11'sd545}},
{{10'sd460, 9'sd-142, 12'sd1917}, {12'sd1940, 11'sd890, 13'sd-2081}, {11'sd934, 13'sd2374, 13'sd-2083}},
{{11'sd1002, 11'sd884, 12'sd-1070}, {13'sd2128, 12'sd-1745, 10'sd457}, {13'sd2128, 12'sd1180, 8'sd109}},
{{13'sd2219, 5'sd-15, 13'sd2316}, {13'sd-2264, 13'sd2370, 12'sd1371}, {11'sd860, 11'sd1021, 12'sd1856}},
{{13'sd2203, 12'sd1915, 11'sd865}, {12'sd1071, 11'sd-992, 10'sd393}, {12'sd-1273, 8'sd126, 12'sd-1774}},
{{10'sd440, 5'sd-11, 10'sd-404}, {12'sd1757, 12'sd1338, 13'sd-3046}, {12'sd-1616, 13'sd-3431, 10'sd352}},
{{13'sd-2816, 12'sd1714, 12'sd1564}, {13'sd2378, 12'sd-1048, 12'sd1821}, {13'sd2619, 13'sd-2609, 13'sd2579}},
{{13'sd-2627, 13'sd2143, 11'sd-740}, {13'sd-2067, 11'sd941, 13'sd-2796}, {11'sd-566, 11'sd872, 13'sd-2637}},
{{11'sd-636, 12'sd-1865, 11'sd967}, {12'sd1356, 13'sd-2188, 13'sd-2227}, {11'sd-938, 10'sd-292, 11'sd-975}},
{{12'sd1494, 11'sd535, 8'sd74}, {11'sd541, 12'sd1946, 13'sd2642}, {10'sd-321, 13'sd2696, 11'sd597}},
{{9'sd-225, 13'sd2285, 12'sd-1806}, {13'sd2578, 12'sd-1274, 12'sd1183}, {12'sd1519, 11'sd-695, 12'sd2014}},
{{13'sd-2219, 11'sd557, 12'sd1346}, {11'sd-873, 12'sd1079, 8'sd-111}, {13'sd2053, 13'sd2080, 12'sd-1674}},
{{11'sd-605, 13'sd-2268, 11'sd-751}, {13'sd2444, 11'sd-866, 10'sd323}, {12'sd1518, 10'sd-420, 10'sd-509}},
{{12'sd-1488, 12'sd-1582, 12'sd1714}, {10'sd439, 12'sd1263, 13'sd2285}, {11'sd-806, 13'sd2077, 13'sd2535}},
{{12'sd-1075, 13'sd2113, 11'sd-881}, {12'sd1474, 12'sd1212, 13'sd2500}, {13'sd2683, 12'sd1937, 12'sd1793}},
{{10'sd407, 9'sd-168, 13'sd2113}, {12'sd1134, 12'sd1818, 12'sd1879}, {13'sd2743, 13'sd2767, 10'sd-356}},
{{13'sd-2878, 12'sd1096, 13'sd2383}, {13'sd2115, 12'sd-1774, 11'sd853}, {12'sd1458, 9'sd167, 12'sd-1307}},
{{13'sd-2459, 12'sd1032, 10'sd-454}, {12'sd1713, 9'sd-255, 12'sd1166}, {13'sd-2086, 12'sd1559, 12'sd1688}},
{{12'sd-1314, 12'sd-1784, 11'sd827}, {9'sd-177, 11'sd660, 12'sd-1900}, {11'sd616, 13'sd-3677, 11'sd763}},
{{12'sd-1068, 13'sd2314, 13'sd-2384}, {11'sd906, 11'sd882, 10'sd399}, {12'sd-1884, 11'sd937, 13'sd-2263}},
{{12'sd-1091, 10'sd463, 9'sd-200}, {11'sd742, 12'sd1324, 13'sd2422}, {13'sd-2395, 12'sd-1209, 10'sd-260}},
{{10'sd370, 12'sd1918, 13'sd-2390}, {12'sd-1153, 13'sd-2161, 13'sd-2343}, {10'sd-374, 12'sd-1891, 11'sd-664}},
{{11'sd-614, 13'sd-2297, 12'sd1220}, {13'sd-2216, 13'sd-2283, 12'sd-1400}, {12'sd1802, 13'sd2343, 12'sd-1329}},
{{8'sd-69, 13'sd2169, 9'sd238}, {9'sd-227, 9'sd175, 13'sd2332}, {13'sd-2545, 12'sd1536, 11'sd666}},
{{9'sd-149, 11'sd573, 11'sd-909}, {13'sd-2437, 12'sd1512, 11'sd-540}, {11'sd-527, 13'sd3223, 13'sd2341}},
{{12'sd1746, 12'sd-1803, 11'sd-654}, {12'sd-1617, 13'sd2193, 11'sd911}, {13'sd2656, 13'sd2588, 13'sd2545}},
{{12'sd-1736, 12'sd-1185, 13'sd-2640}, {13'sd2418, 12'sd-1836, 12'sd-1971}, {13'sd-2338, 13'sd-2713, 12'sd-1331}},
{{13'sd2790, 5'sd10, 13'sd-2064}, {12'sd1300, 11'sd626, 12'sd1958}, {12'sd-1135, 11'sd832, 12'sd-1668}},
{{12'sd-1338, 12'sd-1789, 9'sd-174}, {13'sd-2647, 11'sd-533, 7'sd-36}, {12'sd-1235, 13'sd-2235, 13'sd2139}},
{{11'sd-830, 12'sd-1864, 13'sd-2495}, {13'sd-2620, 13'sd2315, 12'sd1524}, {13'sd-2505, 12'sd2039, 13'sd2401}},
{{13'sd2228, 13'sd-2208, 11'sd622}, {13'sd2192, 13'sd2501, 13'sd-2530}, {13'sd2335, 13'sd-2403, 11'sd-531}},
{{13'sd2540, 9'sd-235, 13'sd-2327}, {13'sd2240, 9'sd152, 12'sd1096}, {12'sd-1562, 10'sd471, 13'sd2951}},
{{13'sd-2454, 10'sd340, 12'sd-1776}, {11'sd-780, 10'sd-373, 12'sd1954}, {12'sd1573, 9'sd-168, 13'sd-2678}},
{{13'sd2186, 12'sd1520, 8'sd-107}, {12'sd1032, 13'sd-2175, 10'sd390}, {12'sd-1885, 13'sd-2777, 12'sd1084}},
{{11'sd756, 12'sd-1865, 13'sd2421}, {11'sd-680, 9'sd-155, 9'sd217}, {10'sd337, 11'sd869, 13'sd2166}},
{{12'sd-1399, 12'sd-1537, 13'sd2489}, {13'sd2081, 13'sd2204, 13'sd-2408}, {12'sd-1580, 13'sd-2277, 10'sd-329}},
{{12'sd2012, 12'sd1800, 11'sd-698}, {12'sd1683, 13'sd2844, 12'sd2007}, {12'sd-1449, 11'sd-838, 12'sd-1898}},
{{11'sd-777, 12'sd1625, 11'sd-771}, {12'sd1308, 13'sd2514, 10'sd-448}, {12'sd-1462, 13'sd-2190, 11'sd555}},
{{12'sd-1935, 13'sd2957, 12'sd2015}, {12'sd1862, 12'sd-1813, 11'sd-884}, {12'sd-1984, 13'sd-2477, 13'sd-3254}},
{{12'sd-1741, 12'sd-1933, 10'sd-508}, {13'sd-2855, 11'sd971, 11'sd720}, {11'sd869, 12'sd-1535, 11'sd889}},
{{13'sd-2831, 12'sd-1174, 12'sd-1862}, {13'sd-2940, 12'sd-1529, 13'sd-2344}, {13'sd-2475, 11'sd-647, 13'sd2303}},
{{12'sd-1424, 12'sd-1717, 13'sd-2673}, {12'sd-1611, 13'sd-2679, 13'sd2312}, {13'sd2091, 6'sd-27, 11'sd912}},
{{11'sd-791, 11'sd-728, 9'sd-228}, {13'sd-2377, 7'sd-62, 12'sd-1942}, {11'sd-655, 12'sd1319, 10'sd383}},
{{12'sd-1554, 13'sd2618, 10'sd345}, {13'sd2667, 12'sd1381, 12'sd1722}, {11'sd-592, 11'sd927, 12'sd-1852}},
{{12'sd-1903, 10'sd456, 12'sd-2023}, {10'sd284, 12'sd-1851, 12'sd-1593}, {8'sd92, 11'sd-628, 12'sd-1733}}},
{
{{13'sd2166, 13'sd2894, 12'sd1951}, {11'sd937, 11'sd904, 11'sd918}, {13'sd-2496, 12'sd1167, 12'sd-1854}},
{{12'sd1920, 13'sd2350, 12'sd1120}, {11'sd-766, 13'sd2288, 12'sd1466}, {10'sd-331, 11'sd-519, 12'sd1243}},
{{12'sd-1263, 11'sd-701, 10'sd-470}, {12'sd-1861, 11'sd768, 9'sd202}, {10'sd-411, 11'sd-842, 13'sd3024}},
{{13'sd2247, 12'sd-1069, 8'sd-126}, {12'sd-1061, 13'sd2251, 11'sd701}, {8'sd-99, 12'sd1392, 10'sd262}},
{{11'sd585, 12'sd-2005, 11'sd996}, {11'sd-747, 12'sd-1316, 12'sd-1485}, {13'sd-2269, 11'sd-889, 13'sd-2191}},
{{13'sd-2589, 12'sd1333, 10'sd400}, {10'sd-299, 13'sd-2105, 12'sd-2027}, {10'sd390, 12'sd1805, 11'sd901}},
{{12'sd-1201, 12'sd-1931, 13'sd2078}, {12'sd1630, 12'sd1308, 9'sd225}, {13'sd2207, 12'sd1553, 13'sd2187}},
{{7'sd51, 12'sd1815, 13'sd-2687}, {8'sd-101, 10'sd486, 13'sd2732}, {12'sd-1194, 10'sd485, 11'sd-644}},
{{11'sd-1016, 10'sd473, 12'sd-1138}, {13'sd-2664, 13'sd-2194, 13'sd2434}, {12'sd-1087, 13'sd-2375, 12'sd-1600}},
{{13'sd-2813, 12'sd-1025, 12'sd-1110}, {12'sd-1892, 10'sd-345, 13'sd-2535}, {3'sd-2, 11'sd545, 11'sd1009}},
{{11'sd599, 8'sd73, 7'sd-56}, {8'sd103, 10'sd-356, 13'sd-2098}, {9'sd-194, 13'sd-2441, 12'sd-1379}},
{{12'sd-1167, 13'sd2442, 11'sd880}, {12'sd1854, 12'sd1514, 13'sd-2413}, {8'sd84, 11'sd-655, 13'sd2081}},
{{12'sd-1118, 10'sd504, 12'sd-1574}, {13'sd-3009, 8'sd-95, 9'sd240}, {11'sd-969, 11'sd-528, 4'sd-7}},
{{12'sd1969, 12'sd-1966, 13'sd2496}, {12'sd1042, 10'sd396, 12'sd-2034}, {11'sd535, 10'sd-505, 13'sd2567}},
{{12'sd-1077, 12'sd1850, 9'sd137}, {10'sd312, 9'sd-177, 7'sd61}, {13'sd2236, 12'sd1975, 12'sd-1067}},
{{11'sd-848, 13'sd3100, 9'sd-140}, {12'sd1894, 12'sd1245, 7'sd43}, {12'sd-1207, 13'sd2396, 11'sd-759}},
{{12'sd-1393, 10'sd373, 4'sd-5}, {8'sd-84, 11'sd702, 13'sd2083}, {12'sd-1047, 11'sd-606, 13'sd-2369}},
{{13'sd-3163, 13'sd-2851, 12'sd1093}, {12'sd-1158, 10'sd344, 13'sd2896}, {13'sd2875, 14'sd4249, 14'sd4720}},
{{10'sd-464, 13'sd-2374, 12'sd1698}, {13'sd-2164, 12'sd1741, 11'sd-1001}, {12'sd-1666, 12'sd-1689, 12'sd1597}},
{{12'sd1512, 13'sd2259, 13'sd2414}, {13'sd-2254, 12'sd-2014, 12'sd1735}, {13'sd2819, 11'sd-1010, 11'sd-584}},
{{11'sd540, 12'sd-1587, 13'sd2778}, {12'sd1730, 10'sd430, 12'sd-1261}, {10'sd498, 13'sd-2609, 13'sd-2067}},
{{10'sd494, 12'sd-1277, 12'sd1792}, {11'sd-999, 13'sd3190, 13'sd-2390}, {13'sd-2512, 13'sd2131, 10'sd271}},
{{13'sd-2119, 12'sd-2036, 11'sd810}, {12'sd1468, 12'sd2038, 12'sd-1225}, {10'sd471, 13'sd-2259, 13'sd-2945}},
{{13'sd2179, 13'sd-2825, 12'sd-1448}, {10'sd-422, 7'sd-58, 12'sd-1402}, {10'sd-260, 13'sd2520, 12'sd-1236}},
{{13'sd-2335, 13'sd-2733, 13'sd2256}, {8'sd117, 9'sd-208, 11'sd-802}, {13'sd-2211, 12'sd2040, 13'sd-2221}},
{{9'sd189, 11'sd951, 12'sd-1948}, {12'sd1496, 13'sd-2497, 10'sd-339}, {13'sd2123, 11'sd-868, 9'sd-157}},
{{12'sd1917, 12'sd1061, 13'sd-2416}, {10'sd-412, 12'sd1612, 12'sd1910}, {12'sd1118, 7'sd44, 11'sd916}},
{{12'sd-1885, 13'sd-2518, 12'sd1700}, {10'sd363, 9'sd-204, 13'sd-2589}, {8'sd117, 12'sd-1116, 13'sd-2479}},
{{11'sd-832, 12'sd-1316, 12'sd-1042}, {12'sd1977, 12'sd1151, 11'sd-1023}, {9'sd-142, 13'sd-2095, 11'sd-1018}},
{{11'sd-616, 11'sd658, 11'sd-879}, {12'sd-1516, 11'sd789, 11'sd774}, {12'sd-1825, 13'sd2296, 12'sd1806}},
{{11'sd518, 9'sd248, 13'sd2271}, {13'sd-2482, 11'sd-551, 10'sd-330}, {12'sd1067, 9'sd-212, 13'sd-2597}},
{{11'sd522, 12'sd-1803, 12'sd-1604}, {11'sd991, 12'sd-1408, 13'sd-2770}, {12'sd1416, 12'sd-1784, 11'sd-917}},
{{11'sd914, 11'sd563, 8'sd85}, {12'sd2013, 13'sd-2782, 9'sd-218}, {13'sd-2472, 11'sd1002, 11'sd583}},
{{12'sd-1552, 11'sd-618, 8'sd-69}, {13'sd-2361, 11'sd925, 11'sd-652}, {13'sd2612, 12'sd1656, 13'sd-2199}},
{{13'sd2162, 11'sd590, 12'sd1297}, {13'sd2866, 12'sd-1274, 11'sd624}, {12'sd-1905, 13'sd2347, 13'sd-2698}},
{{12'sd1268, 12'sd-1474, 12'sd-1254}, {10'sd-485, 13'sd3200, 13'sd2934}, {12'sd1516, 10'sd-261, 10'sd482}},
{{11'sd-925, 13'sd2092, 12'sd-1154}, {12'sd1734, 13'sd-2109, 12'sd-1416}, {13'sd2667, 12'sd-1044, 13'sd2085}},
{{10'sd-377, 13'sd2219, 6'sd-25}, {11'sd953, 12'sd1066, 13'sd-2814}, {9'sd-198, 12'sd-1618, 11'sd-791}},
{{13'sd2278, 7'sd56, 12'sd-1309}, {13'sd2510, 12'sd1759, 12'sd1097}, {13'sd2713, 12'sd2018, 8'sd-84}},
{{11'sd835, 13'sd-2181, 11'sd944}, {13'sd-2434, 12'sd1219, 13'sd-2260}, {11'sd550, 12'sd1250, 7'sd-32}},
{{13'sd-2159, 13'sd2124, 12'sd1542}, {13'sd-3212, 12'sd-1138, 11'sd786}, {11'sd923, 11'sd-735, 11'sd632}},
{{12'sd-1680, 12'sd1274, 12'sd1157}, {12'sd-1513, 12'sd1983, 11'sd713}, {13'sd-2142, 13'sd-2209, 13'sd-2693}},
{{12'sd1361, 7'sd-45, 13'sd-2734}, {10'sd285, 12'sd-1825, 12'sd1064}, {9'sd224, 11'sd577, 11'sd-907}},
{{12'sd-1465, 13'sd2166, 12'sd-1415}, {13'sd2691, 11'sd-512, 8'sd105}, {13'sd2585, 10'sd-328, 11'sd812}},
{{12'sd1194, 12'sd-1417, 11'sd-949}, {10'sd376, 12'sd-1295, 12'sd-1314}, {10'sd-483, 10'sd-482, 13'sd-2493}},
{{13'sd-2518, 13'sd2414, 10'sd357}, {11'sd-598, 10'sd-359, 11'sd-686}, {12'sd-1265, 13'sd-2075, 12'sd-1351}},
{{11'sd-593, 12'sd1524, 12'sd-1323}, {13'sd-2941, 11'sd-858, 12'sd-1057}, {12'sd-1940, 13'sd2673, 13'sd2456}},
{{12'sd-1235, 11'sd-691, 12'sd1805}, {13'sd-2319, 12'sd-1803, 13'sd-2198}, {9'sd203, 13'sd-2699, 13'sd-2255}},
{{12'sd1517, 12'sd1650, 13'sd-2352}, {13'sd2898, 12'sd1582, 12'sd-1651}, {8'sd-124, 12'sd-1698, 10'sd335}},
{{10'sd313, 12'sd1263, 8'sd-82}, {9'sd-193, 12'sd-2045, 12'sd-1443}, {12'sd-1239, 12'sd1414, 8'sd114}},
{{13'sd-2679, 11'sd834, 13'sd-2525}, {13'sd-2194, 13'sd-2265, 13'sd2522}, {7'sd-37, 13'sd2355, 13'sd-3162}},
{{12'sd1785, 10'sd479, 12'sd-1491}, {11'sd843, 12'sd1110, 12'sd1174}, {8'sd-107, 11'sd-869, 11'sd795}},
{{13'sd-2843, 10'sd284, 13'sd2241}, {12'sd-1495, 13'sd-2759, 12'sd1110}, {12'sd-1525, 9'sd165, 13'sd2718}},
{{12'sd-1134, 7'sd-32, 13'sd-2829}, {12'sd-1103, 12'sd-1748, 12'sd-1426}, {9'sd-133, 13'sd-2510, 13'sd-2506}},
{{11'sd-585, 12'sd1284, 13'sd-2663}, {11'sd901, 10'sd367, 6'sd29}, {12'sd1226, 12'sd-1673, 11'sd731}},
{{13'sd-2137, 11'sd-785, 12'sd-1208}, {11'sd-724, 12'sd1076, 11'sd1010}, {11'sd843, 12'sd-1028, 12'sd1269}},
{{12'sd1696, 11'sd650, 12'sd1537}, {13'sd-2747, 11'sd-755, 9'sd139}, {11'sd-996, 11'sd695, 11'sd-606}},
{{12'sd-1285, 12'sd-1193, 7'sd-59}, {12'sd-1571, 7'sd-45, 13'sd-2587}, {11'sd553, 11'sd683, 11'sd601}},
{{12'sd-1973, 13'sd-3642, 13'sd-3026}, {12'sd-1153, 13'sd-2834, 13'sd-3246}, {13'sd2501, 11'sd-912, 13'sd2642}},
{{12'sd1778, 13'sd2760, 10'sd302}, {12'sd-1259, 13'sd2723, 11'sd567}, {13'sd2710, 10'sd455, 13'sd2679}},
{{13'sd-2362, 11'sd648, 10'sd454}, {13'sd-2915, 13'sd2951, 13'sd2074}, {11'sd655, 12'sd1725, 12'sd1289}},
{{9'sd129, 13'sd2825, 13'sd-2296}, {12'sd1121, 13'sd2580, 13'sd-2063}, {12'sd-1034, 11'sd911, 10'sd-287}},
{{13'sd-2267, 12'sd2045, 12'sd1620}, {10'sd-287, 10'sd-511, 12'sd1536}, {13'sd2099, 11'sd536, 10'sd428}},
{{10'sd-430, 12'sd1846, 12'sd1713}, {13'sd2070, 12'sd1059, 11'sd-760}, {12'sd-1519, 12'sd-1456, 12'sd1600}}},
{
{{11'sd584, 12'sd-1173, 12'sd1970}, {12'sd-1569, 9'sd183, 12'sd-1235}, {12'sd1325, 9'sd-232, 7'sd-60}},
{{12'sd1449, 13'sd-2578, 12'sd-1599}, {12'sd-1090, 11'sd557, 11'sd-851}, {11'sd-579, 11'sd876, 13'sd-2648}},
{{11'sd694, 12'sd1509, 12'sd-1151}, {10'sd-441, 12'sd-1107, 11'sd597}, {12'sd1236, 13'sd-2459, 12'sd1100}},
{{13'sd2222, 9'sd-157, 12'sd-1447}, {11'sd829, 10'sd-489, 12'sd1914}, {13'sd2909, 12'sd-1431, 10'sd-258}},
{{13'sd-2299, 9'sd-132, 13'sd-3312}, {13'sd-2077, 10'sd472, 11'sd-871}, {11'sd-799, 11'sd546, 12'sd1402}},
{{13'sd-2314, 9'sd151, 13'sd2164}, {10'sd-416, 12'sd1099, 12'sd1834}, {12'sd-1604, 9'sd148, 11'sd631}},
{{12'sd2008, 12'sd-1775, 13'sd2663}, {11'sd-580, 12'sd-1290, 10'sd422}, {12'sd-1035, 12'sd1358, 12'sd-1642}},
{{13'sd2870, 13'sd2569, 12'sd-1039}, {12'sd1091, 12'sd-1047, 12'sd-1193}, {9'sd-129, 12'sd1850, 13'sd-2240}},
{{10'sd406, 12'sd-1536, 13'sd3190}, {12'sd-1657, 11'sd-1006, 13'sd3286}, {12'sd1989, 13'sd-2501, 7'sd34}},
{{10'sd-399, 10'sd-388, 11'sd540}, {12'sd1161, 11'sd-640, 13'sd3194}, {9'sd-230, 10'sd-385, 12'sd1195}},
{{9'sd189, 12'sd-1458, 13'sd-3913}, {10'sd-376, 10'sd329, 8'sd88}, {13'sd-3270, 14'sd-4197, 14'sd-4764}},
{{12'sd-1704, 13'sd2168, 7'sd39}, {12'sd-1831, 10'sd-401, 12'sd1463}, {10'sd406, 10'sd-385, 12'sd1924}},
{{13'sd2717, 11'sd983, 11'sd-592}, {7'sd38, 12'sd-1893, 11'sd-532}, {12'sd-1833, 13'sd2563, 12'sd2041}},
{{13'sd-2517, 12'sd1435, 12'sd1574}, {11'sd992, 12'sd-1188, 9'sd-207}, {11'sd558, 9'sd-136, 11'sd-962}},
{{12'sd-1332, 13'sd2775, 11'sd-786}, {10'sd-257, 5'sd-14, 12'sd1657}, {13'sd-2590, 12'sd-1194, 12'sd1551}},
{{12'sd-1638, 11'sd-1020, 12'sd-1713}, {11'sd-612, 12'sd-1965, 12'sd1915}, {9'sd-184, 13'sd2461, 12'sd-1597}},
{{13'sd2127, 12'sd-1334, 11'sd-597}, {12'sd1955, 13'sd-3288, 10'sd-374}, {10'sd-492, 12'sd1202, 13'sd-2087}},
{{11'sd-781, 12'sd-1333, 12'sd1623}, {13'sd-2585, 13'sd-2261, 11'sd-731}, {13'sd-2093, 12'sd-1833, 11'sd-675}},
{{13'sd2168, 13'sd2370, 11'sd-775}, {13'sd-2308, 13'sd-2202, 13'sd-2874}, {13'sd2271, 12'sd-1444, 12'sd1342}},
{{11'sd520, 13'sd3458, 11'sd-816}, {11'sd584, 12'sd1323, 11'sd-856}, {13'sd-2471, 12'sd1520, 12'sd-1619}},
{{9'sd131, 13'sd2835, 12'sd1903}, {12'sd-1040, 12'sd1810, 12'sd-1927}, {10'sd-301, 10'sd360, 9'sd184}},
{{13'sd2976, 12'sd-2001, 6'sd-25}, {11'sd-908, 12'sd-1882, 13'sd-2577}, {12'sd1953, 9'sd-202, 9'sd219}},
{{11'sd658, 12'sd1238, 10'sd-489}, {11'sd547, 12'sd1665, 9'sd-155}, {11'sd-668, 10'sd314, 12'sd1320}},
{{12'sd-1073, 13'sd2375, 12'sd-1158}, {11'sd-682, 12'sd-1765, 12'sd1093}, {13'sd2754, 11'sd878, 12'sd-1168}},
{{13'sd-3244, 12'sd-1661, 10'sd-491}, {12'sd1824, 12'sd-1953, 13'sd2128}, {13'sd2713, 13'sd2802, 13'sd3820}},
{{10'sd470, 9'sd-235, 11'sd-703}, {12'sd-1259, 12'sd-1063, 12'sd2025}, {12'sd1661, 13'sd2898, 9'sd149}},
{{10'sd498, 12'sd-1109, 10'sd481}, {11'sd973, 12'sd-1606, 12'sd-1634}, {13'sd2571, 13'sd2614, 12'sd-1531}},
{{11'sd-815, 11'sd-622, 13'sd2060}, {8'sd-82, 9'sd151, 12'sd1584}, {13'sd-2658, 13'sd2490, 10'sd-497}},
{{12'sd1522, 8'sd-107, 12'sd1935}, {12'sd1628, 11'sd-921, 10'sd-456}, {12'sd-1142, 10'sd-391, 10'sd311}},
{{8'sd-109, 12'sd1485, 11'sd638}, {12'sd-1975, 12'sd-1448, 10'sd-464}, {11'sd-789, 12'sd1756, 11'sd550}},
{{11'sd679, 13'sd-2098, 13'sd2216}, {13'sd2499, 9'sd-252, 12'sd1583}, {13'sd-2162, 11'sd-717, 12'sd1555}},
{{12'sd1047, 13'sd-2083, 10'sd-459}, {11'sd916, 12'sd1956, 12'sd1530}, {12'sd-1987, 12'sd-1590, 12'sd-1132}},
{{12'sd-1421, 12'sd1107, 11'sd-562}, {6'sd-24, 12'sd-1038, 13'sd2644}, {13'sd2718, 12'sd1263, 13'sd-2171}},
{{13'sd2071, 13'sd2534, 13'sd2947}, {12'sd1456, 9'sd203, 12'sd1053}, {9'sd-218, 12'sd1966, 13'sd2800}},
{{11'sd672, 12'sd1439, 12'sd-1035}, {12'sd-1466, 12'sd-1555, 12'sd-1701}, {8'sd71, 13'sd2435, 12'sd-1375}},
{{12'sd-1938, 12'sd-2034, 12'sd-1271}, {12'sd-1414, 11'sd-907, 12'sd1460}, {12'sd-1202, 12'sd1989, 12'sd-1463}},
{{11'sd-880, 12'sd-1857, 10'sd-263}, {12'sd-1257, 10'sd-479, 13'sd-2611}, {11'sd684, 8'sd65, 10'sd-331}},
{{13'sd-2792, 9'sd195, 9'sd-164}, {13'sd-2628, 12'sd1124, 10'sd389}, {12'sd-1191, 13'sd-2631, 12'sd-1663}},
{{12'sd-2032, 11'sd-911, 11'sd-702}, {11'sd-996, 12'sd1194, 11'sd-935}, {13'sd-2367, 11'sd-612, 13'sd-2163}},
{{13'sd2583, 13'sd2170, 12'sd-1147}, {13'sd-3181, 13'sd-2385, 6'sd27}, {11'sd-715, 13'sd2225, 12'sd1342}},
{{13'sd2559, 13'sd-2451, 12'sd1834}, {13'sd-2459, 11'sd1011, 7'sd-41}, {11'sd656, 13'sd-2269, 11'sd948}},
{{11'sd907, 13'sd-2515, 12'sd-1343}, {13'sd-2333, 7'sd34, 13'sd-2088}, {12'sd-1994, 11'sd1014, 13'sd2930}},
{{13'sd-2551, 10'sd-416, 12'sd1836}, {9'sd-155, 11'sd-701, 12'sd-1255}, {12'sd-1088, 12'sd1255, 12'sd1102}},
{{10'sd283, 13'sd-2188, 11'sd-809}, {13'sd-2794, 7'sd-51, 12'sd1482}, {10'sd283, 13'sd3287, 12'sd1582}},
{{13'sd2280, 13'sd2165, 13'sd2056}, {12'sd-1493, 12'sd-1737, 12'sd2014}, {12'sd1403, 8'sd75, 12'sd1594}},
{{13'sd-2106, 12'sd-1896, 12'sd-1741}, {10'sd-356, 13'sd2937, 10'sd-380}, {12'sd-1998, 9'sd228, 13'sd2219}},
{{12'sd2017, 11'sd527, 11'sd992}, {13'sd-2253, 11'sd-722, 12'sd-1745}, {13'sd-3191, 9'sd229, 12'sd1501}},
{{11'sd887, 13'sd-2248, 12'sd1645}, {10'sd334, 9'sd208, 12'sd-1754}, {12'sd-1953, 12'sd-1474, 12'sd1853}},
{{13'sd-2196, 8'sd-77, 12'sd-1603}, {13'sd2413, 10'sd300, 11'sd831}, {13'sd2242, 12'sd1852, 12'sd1614}},
{{12'sd1290, 12'sd-1741, 13'sd2133}, {13'sd2531, 9'sd128, 12'sd-1488}, {9'sd171, 9'sd-218, 12'sd-1886}},
{{11'sd-684, 12'sd-1421, 13'sd-2129}, {12'sd1117, 12'sd-1683, 11'sd691}, {9'sd155, 11'sd714, 10'sd302}},
{{8'sd-102, 13'sd-2345, 11'sd-664}, {13'sd2228, 11'sd552, 10'sd-427}, {13'sd2825, 13'sd-2344, 11'sd-726}},
{{11'sd747, 13'sd-3175, 13'sd-2526}, {11'sd-946, 14'sd-4522, 12'sd-1455}, {7'sd40, 14'sd-4304, 13'sd-2095}},
{{9'sd-187, 12'sd-1583, 10'sd-312}, {11'sd-1019, 11'sd845, 11'sd819}, {12'sd-2042, 11'sd-816, 13'sd-2577}},
{{12'sd-1973, 12'sd-1970, 13'sd-2477}, {10'sd267, 12'sd1455, 11'sd-950}, {12'sd-1259, 12'sd1838, 13'sd2190}},
{{13'sd2503, 10'sd352, 13'sd2589}, {12'sd1191, 12'sd1635, 9'sd239}, {13'sd2939, 13'sd-2546, 11'sd-965}},
{{12'sd-1777, 12'sd1766, 13'sd3041}, {12'sd1454, 12'sd-1788, 9'sd138}, {11'sd-860, 12'sd-1811, 9'sd-246}},
{{11'sd-571, 12'sd2040, 5'sd12}, {12'sd1228, 11'sd-810, 12'sd-1326}, {12'sd-1191, 10'sd439, 9'sd-193}},
{{13'sd2280, 13'sd2713, 12'sd-1534}, {11'sd728, 12'sd1952, 10'sd332}, {10'sd-488, 13'sd3156, 11'sd-1009}},
{{9'sd-250, 12'sd-1672, 12'sd1047}, {8'sd-86, 10'sd-360, 3'sd-3}, {12'sd-1629, 11'sd786, 13'sd2980}},
{{11'sd640, 11'sd831, 8'sd121}, {11'sd953, 10'sd-481, 12'sd-1575}, {12'sd-1615, 13'sd2291, 13'sd2461}},
{{11'sd996, 13'sd-2477, 13'sd-2152}, {12'sd-1699, 13'sd-2753, 12'sd-1619}, {12'sd-1184, 12'sd-1465, 10'sd325}},
{{10'sd471, 12'sd-1475, 12'sd1825}, {10'sd-511, 12'sd1567, 13'sd2933}, {10'sd425, 13'sd2639, 11'sd583}},
{{11'sd-867, 11'sd812, 12'sd1564}, {13'sd-2247, 10'sd-405, 12'sd-1042}, {12'sd1593, 12'sd-1450, 13'sd3291}}},
{
{{12'sd1411, 12'sd-1561, 11'sd-1002}, {12'sd1182, 13'sd2191, 12'sd1313}, {13'sd2136, 12'sd-1147, 11'sd-549}},
{{11'sd606, 13'sd-3107, 13'sd3123}, {12'sd-1802, 11'sd-607, 13'sd2201}, {11'sd-994, 14'sd-4417, 12'sd1680}},
{{9'sd170, 13'sd-2838, 13'sd3592}, {13'sd-2074, 12'sd1173, 12'sd-1139}, {11'sd-601, 12'sd-1043, 11'sd-598}},
{{8'sd-95, 11'sd-713, 11'sd864}, {10'sd-312, 13'sd2062, 9'sd198}, {7'sd56, 11'sd674, 12'sd-1119}},
{{8'sd80, 13'sd2656, 12'sd-1218}, {11'sd944, 11'sd-650, 11'sd-691}, {12'sd-1334, 11'sd-905, 11'sd-815}},
{{12'sd1234, 12'sd-1352, 12'sd-1609}, {13'sd-3014, 13'sd2229, 11'sd819}, {12'sd1974, 9'sd132, 11'sd-530}},
{{14'sd4977, 14'sd4908, 13'sd2637}, {13'sd-3766, 10'sd-344, 13'sd-3168}, {10'sd-399, 13'sd-2901, 12'sd-1814}},
{{13'sd4006, 12'sd1997, 13'sd-2409}, {12'sd1479, 12'sd1226, 12'sd-1415}, {9'sd227, 10'sd335, 12'sd1221}},
{{13'sd-3909, 11'sd-828, 13'sd-3201}, {13'sd2890, 13'sd2842, 12'sd1472}, {13'sd4013, 12'sd1508, 13'sd2671}},
{{13'sd3196, 12'sd1994, 13'sd3280}, {12'sd-2010, 13'sd-2611, 11'sd-738}, {13'sd3403, 12'sd1164, 13'sd3429}},
{{13'sd2138, 14'sd5371, 12'sd-1294}, {13'sd3492, 13'sd3987, 12'sd-1071}, {13'sd2678, 9'sd252, 13'sd-3645}},
{{12'sd-1897, 11'sd709, 11'sd638}, {8'sd88, 13'sd-2424, 13'sd-2593}, {11'sd-739, 12'sd2042, 13'sd2101}},
{{12'sd1994, 12'sd1872, 13'sd3964}, {13'sd-2989, 13'sd-2655, 12'sd1986}, {13'sd-3436, 9'sd247, 14'sd4317}},
{{12'sd1208, 12'sd2026, 12'sd-1102}, {11'sd-668, 11'sd775, 9'sd-159}, {13'sd2050, 13'sd2669, 13'sd-2782}},
{{11'sd-852, 12'sd-1797, 12'sd-1897}, {12'sd-1578, 13'sd-2175, 12'sd-1338}, {13'sd-2579, 10'sd-434, 13'sd2084}},
{{11'sd920, 13'sd-2513, 11'sd-744}, {13'sd3418, 12'sd1241, 12'sd-2040}, {12'sd1149, 12'sd-1568, 11'sd609}},
{{12'sd-1608, 12'sd2023, 9'sd-157}, {13'sd2128, 10'sd492, 13'sd2419}, {7'sd49, 11'sd723, 12'sd1556}},
{{10'sd-340, 12'sd1772, 13'sd3865}, {13'sd-3159, 13'sd-3242, 12'sd-1158}, {13'sd-2368, 13'sd-2216, 12'sd-1824}},
{{13'sd3101, 11'sd649, 12'sd-1324}, {12'sd-1974, 13'sd-2323, 13'sd-3036}, {13'sd-2719, 12'sd1205, 12'sd1944}},
{{11'sd-1011, 12'sd1286, 7'sd50}, {12'sd-1935, 11'sd-935, 13'sd3028}, {11'sd-703, 10'sd-301, 12'sd-1596}},
{{12'sd-1204, 13'sd-2593, 12'sd-1616}, {13'sd-2583, 12'sd1965, 10'sd-264}, {12'sd1882, 11'sd845, 12'sd1467}},
{{12'sd1958, 13'sd4021, 12'sd1088}, {11'sd1000, 12'sd1692, 11'sd614}, {12'sd1478, 13'sd-3029, 14'sd-5019}},
{{13'sd2153, 12'sd-1426, 13'sd2194}, {12'sd1263, 9'sd-196, 12'sd-1635}, {10'sd388, 12'sd-1698, 13'sd2288}},
{{11'sd733, 12'sd1638, 12'sd1808}, {10'sd-339, 12'sd-1399, 10'sd-447}, {13'sd2988, 12'sd1599, 13'sd-2394}},
{{13'sd-3100, 13'sd-2636, 13'sd-3062}, {13'sd3402, 13'sd-2590, 13'sd3129}, {12'sd1090, 12'sd2018, 14'sd4713}},
{{13'sd-2061, 13'sd2791, 12'sd-1407}, {13'sd-2565, 12'sd-1097, 11'sd549}, {5'sd-14, 11'sd863, 12'sd-1803}},
{{13'sd-2667, 12'sd-1255, 13'sd-2927}, {12'sd1676, 12'sd1768, 13'sd-2141}, {12'sd1491, 10'sd-396, 10'sd-508}},
{{11'sd702, 12'sd-1354, 12'sd1303}, {11'sd-735, 13'sd-2223, 12'sd1241}, {13'sd2481, 11'sd-833, 12'sd-1669}},
{{11'sd561, 11'sd-591, 13'sd2635}, {11'sd-658, 12'sd-1693, 12'sd1386}, {14'sd-5063, 14'sd-4278, 13'sd-2292}},
{{11'sd-849, 12'sd1389, 12'sd-1494}, {13'sd3634, 13'sd2742, 13'sd-2642}, {12'sd1347, 13'sd2915, 13'sd-2422}},
{{12'sd-1507, 12'sd-1518, 10'sd459}, {12'sd-1955, 11'sd811, 11'sd736}, {11'sd578, 13'sd-2496, 13'sd-2365}},
{{12'sd-1918, 13'sd-3260, 13'sd-2453}, {13'sd-2076, 13'sd-3533, 12'sd-1873}, {12'sd-1484, 14'sd-4449, 13'sd-2763}},
{{13'sd-2414, 13'sd-2311, 12'sd1189}, {13'sd2658, 12'sd-2000, 9'sd-210}, {11'sd-567, 10'sd-483, 13'sd2538}},
{{13'sd-2891, 12'sd1740, 12'sd1605}, {10'sd-340, 6'sd25, 13'sd3165}, {12'sd1381, 12'sd1860, 12'sd1067}},
{{10'sd-507, 12'sd-1212, 9'sd-139}, {11'sd678, 12'sd1563, 11'sd710}, {11'sd-914, 14'sd4140, 11'sd-920}},
{{12'sd-1719, 12'sd1985, 11'sd577}, {11'sd-522, 11'sd-596, 13'sd-2335}, {10'sd-414, 12'sd1636, 13'sd2596}},
{{11'sd-750, 12'sd1288, 13'sd-2343}, {12'sd1478, 13'sd2213, 12'sd1200}, {11'sd-981, 13'sd-2951, 10'sd-312}},
{{13'sd3811, 13'sd-2117, 10'sd256}, {13'sd2466, 9'sd169, 12'sd-2011}, {11'sd709, 13'sd-3594, 12'sd1197}},
{{12'sd-1583, 12'sd1287, 10'sd-446}, {11'sd-792, 13'sd-2996, 5'sd15}, {13'sd-2350, 14'sd-4103, 10'sd359}},
{{13'sd3501, 10'sd-390, 13'sd3674}, {11'sd-601, 13'sd-2479, 13'sd-2835}, {13'sd-2706, 13'sd-3183, 8'sd-122}},
{{13'sd2518, 12'sd-1607, 10'sd488}, {13'sd-2188, 8'sd-112, 10'sd-356}, {12'sd2047, 13'sd-2920, 12'sd1319}},
{{10'sd-290, 10'sd-396, 9'sd-151}, {13'sd2987, 9'sd231, 13'sd-2785}, {13'sd3551, 12'sd2031, 11'sd-778}},
{{10'sd510, 12'sd-1266, 13'sd2076}, {12'sd-1488, 12'sd-1552, 12'sd-1260}, {12'sd1875, 12'sd-1479, 11'sd992}},
{{9'sd-226, 12'sd-1347, 11'sd575}, {11'sd771, 8'sd67, 11'sd-617}, {12'sd-1475, 13'sd2742, 11'sd868}},
{{12'sd-1332, 13'sd2312, 12'sd1687}, {13'sd2655, 13'sd2214, 12'sd-1096}, {12'sd1753, 4'sd5, 13'sd2137}},
{{12'sd1290, 13'sd-2390, 13'sd-2374}, {13'sd3586, 13'sd3059, 9'sd-138}, {13'sd-2511, 13'sd-2835, 13'sd-2683}},
{{13'sd3763, 10'sd-445, 14'sd4127}, {12'sd-1231, 9'sd-206, 11'sd695}, {13'sd-2452, 13'sd-2725, 12'sd-1730}},
{{13'sd2077, 12'sd1462, 13'sd2166}, {12'sd-1358, 12'sd-1751, 13'sd2401}, {11'sd-673, 11'sd613, 9'sd231}},
{{13'sd-2100, 13'sd2364, 10'sd-417}, {12'sd-1225, 13'sd-2088, 13'sd-2077}, {12'sd-1133, 13'sd2165, 12'sd1161}},
{{13'sd3722, 10'sd454, 12'sd1291}, {12'sd1865, 13'sd-2412, 9'sd243}, {12'sd-1574, 13'sd-2227, 8'sd104}},
{{12'sd-1251, 11'sd-850, 13'sd2233}, {13'sd-2979, 13'sd2755, 12'sd1369}, {13'sd-2485, 11'sd957, 13'sd2741}},
{{13'sd-2790, 11'sd-564, 13'sd-3108}, {7'sd-54, 13'sd2713, 12'sd1191}, {10'sd260, 12'sd-1649, 12'sd1251}},
{{14'sd4318, 14'sd4096, 12'sd1251}, {13'sd-2458, 11'sd-921, 11'sd961}, {12'sd-1734, 11'sd-692, 12'sd-1027}},
{{12'sd-1607, 12'sd1194, 13'sd2410}, {13'sd2159, 13'sd-3484, 10'sd341}, {10'sd352, 11'sd-822, 13'sd-2580}},
{{13'sd2630, 11'sd725, 13'sd2468}, {10'sd-413, 12'sd1532, 10'sd-367}, {12'sd1923, 13'sd-2731, 10'sd371}},
{{12'sd-1166, 12'sd-1442, 13'sd2106}, {12'sd-1630, 11'sd-902, 8'sd-120}, {12'sd1839, 12'sd2035, 12'sd-1502}},
{{13'sd-2451, 10'sd-318, 10'sd-485}, {10'sd-272, 11'sd930, 12'sd1575}, {11'sd867, 13'sd-2809, 12'sd1459}},
{{12'sd1303, 13'sd-2682, 12'sd-1241}, {10'sd292, 14'sd-5284, 13'sd-4068}, {12'sd1162, 11'sd967, 13'sd-2176}},
{{10'sd264, 8'sd104, 12'sd-1067}, {12'sd2043, 11'sd971, 13'sd-3375}, {14'sd6419, 13'sd2381, 13'sd2719}},
{{10'sd474, 12'sd-1472, 12'sd1440}, {12'sd-1572, 12'sd1146, 13'sd-2677}, {11'sd604, 11'sd536, 12'sd1092}},
{{12'sd-1736, 11'sd-677, 10'sd-320}, {12'sd-2001, 8'sd67, 13'sd-2485}, {13'sd2080, 10'sd322, 8'sd106}},
{{11'sd-785, 11'sd557, 12'sd-1034}, {7'sd-36, 11'sd1021, 13'sd2250}, {12'sd1099, 13'sd-2182, 10'sd316}},
{{14'sd-5232, 12'sd-1381, 12'sd1498}, {9'sd137, 11'sd-1014, 13'sd3403}, {8'sd-117, 12'sd-1089, 9'sd193}},
{{13'sd-3153, 12'sd1906, 12'sd1341}, {11'sd-604, 11'sd923, 12'sd1790}, {13'sd-2503, 9'sd-139, 13'sd2700}}},
{
{{12'sd-1416, 11'sd706, 13'sd-2073}, {13'sd-2400, 12'sd-1056, 12'sd-1289}, {13'sd-2343, 12'sd-1916, 12'sd-1690}},
{{11'sd-736, 13'sd-2741, 12'sd1040}, {11'sd-716, 13'sd2424, 13'sd2824}, {11'sd884, 10'sd463, 12'sd1461}},
{{13'sd2538, 9'sd137, 9'sd-141}, {12'sd-1414, 13'sd-2587, 10'sd428}, {12'sd1776, 13'sd-3414, 12'sd-1279}},
{{13'sd-2670, 13'sd-2824, 12'sd1123}, {11'sd575, 13'sd2260, 4'sd5}, {11'sd-746, 13'sd2401, 13'sd-2202}},
{{13'sd2431, 11'sd-611, 13'sd-2284}, {11'sd-586, 12'sd-1197, 12'sd1465}, {12'sd-1924, 13'sd-2262, 9'sd-184}},
{{13'sd-2750, 10'sd269, 11'sd-764}, {12'sd2039, 12'sd1648, 13'sd2401}, {13'sd2104, 13'sd-2364, 8'sd-111}},
{{13'sd2329, 13'sd2366, 12'sd-1626}, {13'sd-2517, 12'sd-1995, 11'sd-738}, {10'sd327, 12'sd-1738, 13'sd-2205}},
{{12'sd1624, 11'sd-891, 11'sd822}, {11'sd616, 13'sd-2535, 12'sd1223}, {13'sd2996, 11'sd-692, 13'sd-2490}},
{{10'sd-414, 13'sd-2676, 12'sd1568}, {12'sd-1884, 13'sd2349, 13'sd-2712}, {12'sd1662, 11'sd1001, 13'sd-2737}},
{{12'sd-1798, 12'sd-2010, 12'sd-1106}, {11'sd742, 11'sd818, 9'sd-142}, {11'sd642, 12'sd1643, 13'sd2329}},
{{13'sd2587, 12'sd-1309, 10'sd-463}, {12'sd1317, 10'sd-410, 13'sd2081}, {11'sd-666, 12'sd1931, 6'sd-20}},
{{11'sd597, 11'sd794, 12'sd-1263}, {13'sd-2283, 11'sd600, 9'sd243}, {10'sd499, 13'sd2727, 12'sd1899}},
{{9'sd-133, 12'sd1704, 12'sd-1227}, {12'sd-1588, 12'sd-1579, 12'sd-1029}, {12'sd1946, 12'sd1645, 13'sd2748}},
{{11'sd-913, 10'sd-378, 11'sd-940}, {13'sd-2591, 12'sd-1877, 12'sd-1967}, {13'sd2471, 13'sd-2558, 12'sd1566}},
{{13'sd-2638, 13'sd-2667, 10'sd321}, {12'sd1156, 10'sd-493, 10'sd450}, {12'sd1727, 10'sd-386, 10'sd-358}},
{{9'sd161, 10'sd289, 12'sd-1322}, {12'sd1401, 12'sd-1486, 12'sd-1395}, {7'sd52, 12'sd-1139, 13'sd2215}},
{{13'sd-2088, 10'sd-298, 13'sd-2200}, {12'sd-1471, 11'sd759, 12'sd-1112}, {11'sd-867, 13'sd2347, 10'sd-416}},
{{10'sd-331, 10'sd-403, 11'sd786}, {12'sd1162, 13'sd-2199, 9'sd196}, {12'sd-1372, 13'sd-2088, 12'sd1102}},
{{12'sd1909, 12'sd1283, 12'sd1825}, {12'sd-1123, 13'sd2525, 12'sd-1288}, {10'sd-476, 11'sd-745, 11'sd-708}},
{{12'sd1594, 11'sd-575, 12'sd-1188}, {8'sd125, 12'sd1806, 12'sd-2045}, {12'sd1933, 11'sd624, 12'sd1497}},
{{12'sd-1987, 13'sd-2572, 12'sd-1400}, {13'sd2491, 12'sd-1464, 13'sd-2658}, {13'sd2447, 12'sd-1080, 4'sd-7}},
{{11'sd-662, 12'sd1193, 12'sd-1219}, {11'sd-691, 13'sd2434, 12'sd1250}, {12'sd1137, 11'sd589, 13'sd2556}},
{{10'sd-350, 13'sd2256, 13'sd2288}, {13'sd-2443, 13'sd-2210, 12'sd1446}, {11'sd1009, 12'sd-1263, 11'sd-822}},
{{9'sd-206, 13'sd-2460, 11'sd969}, {12'sd1113, 11'sd692, 10'sd-258}, {12'sd1411, 12'sd1710, 10'sd395}},
{{13'sd-2470, 13'sd2176, 10'sd488}, {11'sd-892, 12'sd2008, 13'sd2704}, {11'sd918, 9'sd179, 11'sd798}},
{{8'sd-91, 13'sd-2621, 10'sd-462}, {5'sd14, 12'sd1753, 9'sd-157}, {13'sd2699, 13'sd-2090, 12'sd-1426}},
{{12'sd1106, 12'sd-1881, 12'sd-1842}, {12'sd-1640, 9'sd248, 11'sd-1009}, {13'sd2614, 12'sd-1851, 12'sd-1885}},
{{13'sd2749, 12'sd-1554, 13'sd-2415}, {11'sd940, 11'sd746, 9'sd-239}, {13'sd-2155, 11'sd1009, 11'sd607}},
{{11'sd604, 9'sd-167, 13'sd-2477}, {10'sd-270, 12'sd-1257, 13'sd-2673}, {11'sd704, 12'sd-1518, 13'sd2542}},
{{12'sd-1177, 11'sd-769, 13'sd2427}, {10'sd314, 13'sd2335, 13'sd2282}, {10'sd-505, 13'sd2306, 13'sd2590}},
{{12'sd-1969, 12'sd-1216, 13'sd2229}, {12'sd-1852, 12'sd1143, 11'sd-868}, {9'sd-159, 13'sd2674, 13'sd2113}},
{{12'sd-1491, 13'sd2497, 10'sd258}, {11'sd828, 12'sd1476, 13'sd2288}, {9'sd-234, 12'sd-1572, 13'sd-2476}},
{{11'sd-1017, 13'sd2478, 13'sd-2680}, {12'sd-1971, 13'sd-2423, 12'sd1388}, {13'sd2515, 13'sd-2060, 12'sd-1360}},
{{12'sd-1547, 12'sd-1068, 13'sd2453}, {13'sd2558, 12'sd1913, 11'sd772}, {12'sd-1041, 13'sd-2316, 13'sd-2736}},
{{11'sd-1017, 12'sd1461, 12'sd-1908}, {13'sd2434, 13'sd-2134, 12'sd1837}, {11'sd535, 12'sd-2005, 12'sd1388}},
{{13'sd2420, 12'sd1096, 11'sd760}, {13'sd2153, 12'sd-1036, 12'sd2004}, {11'sd-1001, 10'sd441, 12'sd1385}},
{{12'sd-1595, 13'sd-2856, 11'sd-604}, {13'sd-2122, 12'sd1626, 12'sd1087}, {11'sd965, 6'sd-28, 10'sd492}},
{{11'sd584, 11'sd-948, 11'sd893}, {9'sd-235, 12'sd1668, 12'sd-1230}, {12'sd1934, 12'sd-1132, 11'sd-590}},
{{13'sd-2911, 13'sd3015, 12'sd-1930}, {12'sd1400, 12'sd1984, 13'sd2655}, {12'sd-1977, 12'sd1561, 12'sd-1622}},
{{13'sd-2246, 12'sd1164, 9'sd188}, {13'sd-2224, 11'sd818, 12'sd-1034}, {13'sd-2457, 12'sd1398, 12'sd-1829}},
{{10'sd326, 11'sd-556, 11'sd906}, {13'sd2769, 13'sd-2453, 12'sd-1849}, {11'sd948, 10'sd389, 11'sd-714}},
{{11'sd-816, 12'sd1819, 12'sd1047}, {11'sd850, 13'sd2710, 10'sd501}, {10'sd-258, 13'sd-2313, 13'sd-2462}},
{{10'sd296, 12'sd1416, 12'sd-2015}, {12'sd1116, 12'sd-1897, 11'sd557}, {12'sd-1529, 11'sd-622, 11'sd758}},
{{13'sd-2811, 10'sd348, 13'sd-2459}, {12'sd-2011, 13'sd2680, 12'sd1368}, {12'sd1407, 13'sd2330, 12'sd-1187}},
{{12'sd-1910, 12'sd-1640, 12'sd1486}, {13'sd2154, 11'sd-529, 8'sd-126}, {10'sd339, 12'sd1610, 13'sd-2513}},
{{12'sd-1558, 12'sd-1088, 12'sd-1692}, {11'sd-929, 13'sd-2691, 12'sd-1659}, {9'sd169, 12'sd1229, 12'sd1326}},
{{9'sd-250, 10'sd-436, 12'sd-1493}, {11'sd-520, 13'sd-2436, 12'sd1188}, {12'sd1650, 11'sd808, 13'sd2166}},
{{11'sd-872, 12'sd1631, 9'sd-252}, {12'sd-1189, 13'sd-2382, 8'sd123}, {3'sd-3, 13'sd-2358, 11'sd-767}},
{{13'sd-2575, 12'sd1570, 11'sd657}, {13'sd2313, 12'sd1532, 8'sd113}, {10'sd-325, 12'sd1556, 12'sd-1736}},
{{11'sd973, 12'sd1408, 11'sd-573}, {13'sd-2105, 12'sd-1800, 11'sd878}, {10'sd260, 13'sd-2467, 13'sd2281}},
{{12'sd-1118, 11'sd743, 13'sd-2617}, {12'sd1405, 12'sd-1862, 12'sd1070}, {13'sd2433, 9'sd234, 13'sd2056}},
{{11'sd-968, 13'sd-2706, 10'sd-390}, {12'sd1102, 12'sd-1103, 10'sd-385}, {12'sd-1957, 13'sd-2275, 11'sd697}},
{{13'sd2129, 12'sd1393, 12'sd1544}, {11'sd526, 12'sd1979, 11'sd-698}, {13'sd-2867, 11'sd578, 9'sd239}},
{{11'sd-1011, 13'sd-2164, 12'sd1519}, {11'sd-767, 12'sd1300, 12'sd1320}, {12'sd1530, 12'sd-1432, 13'sd2135}},
{{13'sd2443, 10'sd-309, 13'sd2328}, {13'sd2048, 11'sd-707, 12'sd-1760}, {12'sd-1891, 13'sd2361, 10'sd290}},
{{10'sd-485, 12'sd1374, 10'sd-349}, {12'sd1557, 10'sd-345, 10'sd491}, {13'sd-2287, 9'sd152, 13'sd-2706}},
{{11'sd-715, 12'sd-1098, 7'sd62}, {12'sd1742, 12'sd-1254, 12'sd-1530}, {12'sd-1075, 12'sd1132, 11'sd993}},
{{13'sd3765, 11'sd552, 8'sd-69}, {12'sd-1991, 11'sd-534, 10'sd-470}, {13'sd-3336, 12'sd1813, 7'sd-47}},
{{13'sd3384, 12'sd1101, 12'sd-1977}, {11'sd959, 12'sd-1037, 12'sd2019}, {13'sd2544, 12'sd-1733, 12'sd1345}},
{{13'sd-2561, 12'sd-1526, 12'sd1428}, {12'sd-1828, 12'sd1437, 13'sd2640}, {11'sd-862, 9'sd-167, 12'sd1582}},
{{11'sd-614, 10'sd478, 11'sd-588}, {11'sd808, 12'sd-1867, 10'sd-306}, {12'sd1364, 11'sd-968, 13'sd3024}},
{{7'sd-38, 10'sd-272, 11'sd928}, {13'sd2136, 12'sd1802, 10'sd-341}, {13'sd2105, 12'sd-1510, 13'sd2609}},
{{11'sd-869, 10'sd478, 12'sd1046}, {12'sd1110, 10'sd-316, 8'sd103}, {12'sd-1757, 11'sd651, 13'sd-2196}},
{{6'sd-16, 13'sd2500, 12'sd-1272}, {12'sd-1274, 12'sd-1199, 12'sd-1607}, {12'sd-1275, 13'sd2643, 9'sd195}}},
{
{{12'sd-1657, 11'sd972, 11'sd881}, {13'sd2140, 12'sd1518, 10'sd-404}, {13'sd2360, 11'sd-563, 11'sd700}},
{{13'sd-2963, 13'sd-2159, 11'sd932}, {11'sd-563, 11'sd639, 10'sd359}, {10'sd293, 10'sd-265, 12'sd2022}},
{{13'sd-3467, 13'sd-2875, 10'sd304}, {13'sd-2169, 11'sd-1021, 11'sd-681}, {13'sd3378, 11'sd981, 10'sd420}},
{{12'sd-2002, 12'sd1703, 13'sd-2922}, {12'sd1179, 12'sd-1612, 11'sd-923}, {8'sd115, 7'sd55, 12'sd-1163}},
{{7'sd-33, 13'sd-2449, 10'sd-284}, {13'sd-3080, 13'sd-3247, 13'sd-3269}, {11'sd-854, 13'sd-2798, 12'sd1306}},
{{13'sd2545, 11'sd604, 12'sd1689}, {13'sd-2694, 9'sd-131, 11'sd-521}, {11'sd774, 12'sd1466, 12'sd-1369}},
{{12'sd-1360, 12'sd1239, 13'sd2050}, {11'sd1001, 11'sd592, 13'sd3879}, {12'sd1272, 12'sd-1475, 11'sd942}},
{{12'sd-1904, 12'sd1712, 13'sd-2811}, {13'sd-3444, 13'sd-2094, 13'sd-2323}, {12'sd1363, 12'sd1193, 9'sd-213}},
{{13'sd2873, 13'sd-2566, 9'sd233}, {9'sd-185, 12'sd1296, 11'sd-1009}, {12'sd1643, 12'sd-1661, 11'sd-754}},
{{12'sd1149, 12'sd-1693, 12'sd1264}, {13'sd2193, 12'sd1486, 10'sd-409}, {13'sd3699, 12'sd-1909, 13'sd3779}},
{{13'sd4078, 12'sd-1903, 13'sd3273}, {8'sd78, 13'sd-2682, 13'sd-2224}, {13'sd-2704, 14'sd-6173, 14'sd-4681}},
{{13'sd2590, 10'sd368, 12'sd1474}, {13'sd-2718, 12'sd-1545, 11'sd559}, {11'sd-557, 12'sd2033, 13'sd-3172}},
{{14'sd4154, 13'sd2899, 13'sd2255}, {6'sd26, 10'sd427, 10'sd431}, {12'sd1625, 12'sd1266, 10'sd-279}},
{{12'sd-1454, 12'sd1752, 12'sd1196}, {12'sd-1926, 12'sd1198, 13'sd-3081}, {12'sd-1841, 13'sd-2279, 12'sd-1307}},
{{13'sd-2639, 13'sd-2972, 13'sd2691}, {12'sd1175, 12'sd1447, 12'sd1823}, {12'sd-1565, 10'sd-362, 12'sd1522}},
{{13'sd-2144, 12'sd-1419, 10'sd448}, {13'sd-2293, 12'sd-1686, 13'sd-2187}, {11'sd667, 11'sd948, 12'sd-1832}},
{{13'sd2834, 5'sd10, 13'sd-2231}, {10'sd444, 10'sd-501, 13'sd3089}, {11'sd-1006, 12'sd1552, 13'sd2746}},
{{13'sd-3040, 12'sd-1753, 13'sd-2146}, {12'sd1399, 12'sd2030, 13'sd3527}, {14'sd4836, 9'sd-159, 13'sd3207}},
{{11'sd923, 11'sd634, 9'sd232}, {11'sd-631, 12'sd1382, 12'sd1904}, {12'sd-1974, 10'sd-337, 10'sd-283}},
{{8'sd-71, 7'sd-62, 13'sd-3413}, {12'sd-1215, 12'sd1434, 9'sd212}, {12'sd1047, 10'sd292, 12'sd-1671}},
{{12'sd-1209, 13'sd-2876, 10'sd-500}, {11'sd-765, 11'sd-703, 11'sd-930}, {13'sd2227, 11'sd-548, 12'sd-1500}},
{{11'sd861, 9'sd178, 10'sd303}, {10'sd-382, 13'sd-2194, 12'sd1787}, {11'sd-658, 13'sd-2219, 12'sd-1858}},
{{12'sd-1439, 10'sd480, 9'sd235}, {12'sd-1656, 12'sd1250, 11'sd941}, {11'sd-1002, 10'sd457, 12'sd-1439}},
{{12'sd1199, 12'sd-1171, 13'sd-2077}, {13'sd2343, 12'sd-1636, 12'sd2026}, {12'sd-1074, 11'sd600, 12'sd-1086}},
{{12'sd-1528, 12'sd-1092, 13'sd3068}, {13'sd2176, 11'sd-813, 12'sd1357}, {12'sd1233, 13'sd2737, 12'sd1451}},
{{9'sd219, 12'sd1937, 12'sd-1296}, {12'sd1681, 13'sd-2655, 12'sd1805}, {13'sd-2529, 13'sd2125, 12'sd-1351}},
{{11'sd552, 8'sd-84, 12'sd1119}, {13'sd2435, 13'sd-2378, 12'sd1048}, {13'sd2579, 11'sd-619, 13'sd-3521}},
{{11'sd-725, 12'sd1702, 13'sd-3023}, {12'sd-1759, 12'sd1991, 11'sd872}, {10'sd399, 8'sd90, 13'sd-2633}},
{{13'sd3048, 12'sd2017, 13'sd-2977}, {12'sd-1892, 12'sd1316, 11'sd954}, {13'sd-2369, 10'sd-380, 12'sd2011}},
{{10'sd325, 12'sd-1635, 13'sd-2144}, {13'sd2095, 13'sd2980, 12'sd-1750}, {13'sd-3083, 13'sd-2127, 13'sd-2755}},
{{13'sd2700, 12'sd1317, 11'sd558}, {13'sd2109, 13'sd-2848, 12'sd-1283}, {13'sd2072, 12'sd1937, 13'sd2409}},
{{13'sd-2838, 11'sd-654, 14'sd-4787}, {11'sd576, 10'sd416, 13'sd-2125}, {12'sd-1894, 13'sd-2294, 12'sd-1971}},
{{11'sd803, 13'sd-2146, 12'sd1687}, {13'sd-2445, 7'sd-50, 13'sd2176}, {12'sd1078, 8'sd-100, 13'sd3572}},
{{12'sd1647, 11'sd640, 10'sd-324}, {11'sd792, 12'sd-1123, 11'sd-847}, {13'sd-2339, 13'sd2511, 9'sd171}},
{{11'sd-709, 12'sd-1144, 12'sd1377}, {12'sd-1858, 12'sd-1657, 11'sd-972}, {13'sd-2236, 13'sd2631, 12'sd-1504}},
{{13'sd2810, 11'sd924, 12'sd-1969}, {11'sd816, 13'sd-2322, 13'sd-2369}, {12'sd1146, 9'sd-140, 13'sd-2884}},
{{8'sd92, 13'sd-3356, 13'sd-2175}, {13'sd-2634, 13'sd-2965, 13'sd-2718}, {13'sd2062, 13'sd-2330, 11'sd564}},
{{13'sd-2289, 11'sd805, 13'sd2271}, {13'sd-3342, 13'sd3735, 11'sd-552}, {13'sd-3621, 11'sd735, 12'sd-1335}},
{{12'sd-1226, 13'sd-2563, 12'sd-1291}, {13'sd-3016, 12'sd-1428, 12'sd-1062}, {12'sd-1103, 14'sd-5024, 12'sd-1186}},
{{13'sd2667, 12'sd1541, 13'sd2118}, {11'sd972, 12'sd-1208, 10'sd-370}, {13'sd-3342, 12'sd-1890, 13'sd2576}},
{{12'sd-1396, 13'sd-2321, 9'sd134}, {12'sd1450, 12'sd-2033, 13'sd2411}, {12'sd-1448, 10'sd504, 11'sd-514}},
{{12'sd-1927, 12'sd-1799, 11'sd-558}, {13'sd2149, 10'sd418, 13'sd2483}, {11'sd1014, 12'sd1510, 12'sd-1545}},
{{13'sd-2797, 13'sd2061, 12'sd1766}, {12'sd-1210, 12'sd-1960, 13'sd-2078}, {12'sd-1815, 10'sd424, 13'sd-3790}},
{{13'sd3693, 12'sd-1760, 11'sd-926}, {12'sd-1201, 12'sd1029, 14'sd-4958}, {12'sd-1053, 14'sd-4764, 14'sd-5492}},
{{12'sd-1942, 11'sd689, 13'sd3132}, {13'sd2108, 13'sd2281, 8'sd69}, {13'sd-2070, 12'sd-1273, 10'sd434}},
{{9'sd-237, 12'sd1301, 10'sd310}, {11'sd-905, 12'sd-1809, 13'sd-2571}, {11'sd-732, 10'sd-281, 6'sd25}},
{{11'sd-841, 12'sd-1803, 13'sd-2168}, {11'sd-707, 12'sd1083, 12'sd1948}, {11'sd731, 12'sd-1131, 13'sd2200}},
{{12'sd-1280, 11'sd-528, 12'sd-1331}, {11'sd794, 10'sd-324, 13'sd2103}, {13'sd2319, 13'sd2418, 13'sd-2134}},
{{11'sd-979, 13'sd2345, 7'sd45}, {12'sd-1608, 10'sd-410, 12'sd1372}, {12'sd1544, 11'sd-747, 13'sd-2122}},
{{13'sd2476, 12'sd-1569, 13'sd2867}, {12'sd1949, 10'sd364, 10'sd406}, {12'sd1513, 13'sd2857, 13'sd2866}},
{{9'sd214, 13'sd2891, 12'sd1982}, {11'sd-777, 12'sd-1870, 13'sd-2438}, {13'sd2106, 12'sd-2021, 9'sd-136}},
{{13'sd2584, 10'sd-393, 13'sd2056}, {9'sd144, 11'sd819, 12'sd1610}, {13'sd2471, 12'sd1726, 11'sd-952}},
{{13'sd-3071, 13'sd3073, 9'sd217}, {7'sd-46, 8'sd-93, 10'sd-302}, {12'sd-1966, 12'sd1902, 13'sd3172}},
{{13'sd-2810, 13'sd-2868, 13'sd-2415}, {11'sd-675, 12'sd1038, 13'sd2453}, {13'sd2692, 11'sd-851, 9'sd-198}},
{{13'sd-2209, 13'sd-2337, 10'sd280}, {11'sd738, 10'sd343, 13'sd2242}, {9'sd-175, 13'sd-2154, 9'sd185}},
{{12'sd1816, 12'sd-2045, 13'sd2678}, {8'sd-122, 7'sd-50, 13'sd3213}, {13'sd2570, 13'sd2190, 4'sd6}},
{{12'sd1867, 10'sd-260, 9'sd239}, {13'sd-3658, 13'sd-3151, 12'sd1050}, {11'sd629, 13'sd3330, 9'sd-173}},
{{12'sd-1956, 13'sd2455, 12'sd1439}, {10'sd-472, 11'sd-755, 13'sd2185}, {12'sd1417, 11'sd559, 12'sd1958}},
{{13'sd3231, 10'sd443, 12'sd-1230}, {12'sd1075, 13'sd2197, 11'sd750}, {11'sd-1022, 13'sd2757, 12'sd-1980}},
{{12'sd-1930, 12'sd1532, 12'sd-1757}, {8'sd81, 13'sd2190, 12'sd1799}, {10'sd-346, 7'sd62, 13'sd-2386}},
{{13'sd-2753, 13'sd-2075, 11'sd-888}, {11'sd767, 11'sd888, 12'sd-1592}, {12'sd1458, 11'sd-733, 10'sd-452}},
{{11'sd863, 12'sd1709, 13'sd2156}, {12'sd1166, 12'sd1683, 11'sd-598}, {12'sd-1151, 12'sd1090, 12'sd-1833}},
{{12'sd1923, 12'sd-1308, 12'sd1686}, {12'sd1300, 11'sd-530, 12'sd-1502}, {12'sd1151, 13'sd2250, 12'sd-1311}},
{{12'sd2013, 12'sd-1304, 11'sd969}, {12'sd-1093, 13'sd2060, 10'sd-452}, {11'sd770, 10'sd466, 13'sd2736}}},
{
{{12'sd1936, 12'sd2046, 9'sd199}, {12'sd1538, 10'sd-349, 13'sd2814}, {12'sd1179, 12'sd1637, 12'sd-1424}},
{{13'sd-2986, 13'sd-2522, 12'sd-1226}, {10'sd320, 11'sd-526, 12'sd-1377}, {13'sd-2343, 12'sd1512, 10'sd-430}},
{{13'sd-3761, 11'sd-636, 13'sd-2602}, {13'sd2905, 13'sd3131, 11'sd643}, {12'sd1427, 12'sd1573, 12'sd1238}},
{{9'sd-229, 10'sd-310, 12'sd1568}, {11'sd-606, 9'sd-139, 12'sd-1890}, {12'sd1427, 12'sd1354, 12'sd1941}},
{{12'sd-1416, 11'sd-797, 12'sd1340}, {10'sd-411, 11'sd-787, 11'sd-588}, {13'sd-2405, 12'sd-1255, 12'sd-1999}},
{{13'sd-2107, 12'sd-1509, 11'sd-928}, {9'sd230, 13'sd-2638, 11'sd549}, {11'sd718, 9'sd-142, 8'sd-125}},
{{11'sd-828, 11'sd-844, 12'sd-1710}, {13'sd-2206, 11'sd-842, 8'sd-69}, {12'sd1684, 11'sd-678, 12'sd1035}},
{{13'sd-2435, 12'sd1688, 13'sd-2660}, {13'sd-2462, 10'sd-386, 10'sd511}, {11'sd-775, 12'sd1625, 11'sd641}},
{{12'sd-1981, 13'sd-2307, 10'sd468}, {12'sd1318, 9'sd221, 12'sd1792}, {11'sd669, 13'sd3166, 12'sd2029}},
{{10'sd267, 10'sd-308, 8'sd-92}, {13'sd2118, 12'sd1337, 13'sd-2302}, {11'sd-699, 12'sd1637, 12'sd1687}},
{{14'sd4831, 11'sd758, 13'sd2067}, {13'sd3469, 13'sd-2735, 10'sd369}, {13'sd2707, 12'sd-1428, 13'sd3844}},
{{10'sd413, 13'sd2540, 10'sd-480}, {13'sd2340, 11'sd858, 10'sd467}, {12'sd-1818, 12'sd-1903, 12'sd-1202}},
{{12'sd-1159, 11'sd896, 13'sd-2628}, {10'sd350, 11'sd551, 12'sd-1647}, {12'sd-1845, 11'sd-690, 13'sd2318}},
{{12'sd1350, 13'sd-2137, 12'sd-1144}, {13'sd-2727, 13'sd2478, 12'sd-1086}, {13'sd-2168, 11'sd-909, 13'sd-2062}},
{{13'sd3461, 6'sd21, 12'sd1065}, {11'sd951, 13'sd-2408, 13'sd-2314}, {9'sd234, 12'sd-1183, 11'sd912}},
{{12'sd1872, 12'sd1884, 11'sd-974}, {12'sd1569, 11'sd533, 12'sd-1228}, {12'sd1628, 13'sd-2118, 13'sd-2601}},
{{13'sd-2839, 11'sd635, 13'sd2104}, {13'sd-2157, 12'sd-1209, 13'sd-2400}, {10'sd-266, 12'sd1811, 13'sd-2306}},
{{8'sd-75, 12'sd1278, 12'sd1436}, {11'sd926, 7'sd57, 11'sd1012}, {13'sd2497, 13'sd3225, 13'sd3901}},
{{11'sd516, 13'sd2416, 11'sd514}, {12'sd1346, 12'sd1740, 12'sd-1719}, {12'sd-1622, 10'sd278, 11'sd-521}},
{{13'sd2212, 12'sd1558, 8'sd77}, {12'sd1075, 12'sd1658, 10'sd496}, {10'sd326, 12'sd-1993, 10'sd469}},
{{10'sd-473, 11'sd1010, 11'sd-798}, {12'sd-1965, 12'sd-1720, 13'sd-2181}, {9'sd-153, 12'sd1836, 12'sd-1603}},
{{7'sd-52, 11'sd693, 9'sd232}, {12'sd-1779, 13'sd-3039, 9'sd-155}, {12'sd-1492, 13'sd-3599, 13'sd-2206}},
{{11'sd-631, 8'sd-99, 12'sd1619}, {13'sd3057, 12'sd-1137, 13'sd-2111}, {12'sd-1483, 11'sd-674, 12'sd-1520}},
{{12'sd1288, 8'sd71, 12'sd-1881}, {12'sd-1540, 12'sd-1922, 13'sd2439}, {12'sd1585, 13'sd2676, 12'sd-1184}},
{{12'sd1608, 10'sd329, 10'sd448}, {11'sd641, 10'sd-311, 9'sd-133}, {12'sd-1700, 10'sd-364, 11'sd-599}},
{{13'sd2577, 11'sd969, 13'sd-2056}, {6'sd-28, 11'sd548, 12'sd1054}, {13'sd-2255, 13'sd-2430, 12'sd-2002}},
{{12'sd1089, 10'sd-298, 11'sd-556}, {12'sd-1616, 12'sd1952, 13'sd2124}, {12'sd-1308, 11'sd717, 12'sd-1465}},
{{13'sd-2187, 12'sd-1421, 9'sd167}, {13'sd-2333, 12'sd-1732, 7'sd-51}, {13'sd-2662, 11'sd605, 12'sd2004}},
{{12'sd-1665, 12'sd-1127, 13'sd-2982}, {11'sd791, 12'sd1848, 9'sd249}, {13'sd2708, 12'sd1738, 12'sd1628}},
{{11'sd700, 13'sd-2817, 10'sd-304}, {12'sd-1480, 13'sd2802, 11'sd-758}, {13'sd-2843, 13'sd-2887, 13'sd-3294}},
{{12'sd1960, 11'sd-934, 12'sd-1926}, {12'sd-1299, 13'sd-2739, 8'sd-101}, {12'sd-1961, 12'sd-1312, 8'sd72}},
{{12'sd-1027, 12'sd1919, 12'sd1690}, {12'sd-1866, 11'sd-774, 10'sd-308}, {9'sd150, 13'sd2778, 12'sd1712}},
{{12'sd-1052, 13'sd2763, 11'sd662}, {13'sd2570, 12'sd-1343, 11'sd-673}, {12'sd1926, 12'sd1840, 12'sd1971}},
{{9'sd-177, 12'sd1775, 10'sd-408}, {12'sd-1882, 13'sd2206, 13'sd2199}, {12'sd-1301, 12'sd2025, 13'sd2391}},
{{12'sd1546, 11'sd964, 12'sd1973}, {10'sd-326, 10'sd428, 12'sd-1765}, {12'sd1859, 13'sd-2609, 13'sd-2976}},
{{12'sd-1513, 12'sd-1428, 12'sd1813}, {13'sd-2075, 11'sd-791, 13'sd2571}, {10'sd-307, 10'sd-327, 11'sd513}},
{{13'sd-2311, 12'sd-1810, 12'sd-1898}, {12'sd1589, 12'sd1137, 9'sd-160}, {12'sd1185, 11'sd-679, 12'sd-1623}},
{{9'sd184, 9'sd228, 11'sd547}, {11'sd572, 13'sd2172, 12'sd-2000}, {12'sd1597, 11'sd-853, 13'sd2262}},
{{12'sd1968, 6'sd-20, 12'sd-1032}, {12'sd1364, 13'sd-2676, 13'sd2141}, {11'sd-731, 13'sd2973, 11'sd567}},
{{10'sd495, 7'sd47, 12'sd-1489}, {13'sd-2605, 9'sd-243, 10'sd459}, {13'sd2794, 12'sd1051, 13'sd2852}},
{{12'sd1842, 13'sd2607, 12'sd1310}, {9'sd-245, 12'sd1701, 12'sd1274}, {12'sd1467, 11'sd745, 12'sd-1582}},
{{12'sd-1546, 13'sd2190, 13'sd2209}, {12'sd1558, 12'sd2013, 12'sd-1392}, {6'sd30, 13'sd2269, 13'sd2433}},
{{13'sd2422, 11'sd-780, 13'sd-2755}, {12'sd-1615, 12'sd1466, 10'sd-348}, {13'sd-2322, 11'sd975, 12'sd1229}},
{{11'sd-846, 11'sd-587, 11'sd-560}, {13'sd-2907, 11'sd-577, 12'sd-1912}, {12'sd-1188, 11'sd774, 5'sd-15}},
{{9'sd158, 12'sd1046, 11'sd-816}, {12'sd1413, 13'sd2396, 11'sd-779}, {13'sd3186, 8'sd-108, 12'sd-1724}},
{{12'sd-1684, 12'sd-1620, 11'sd-532}, {12'sd1369, 12'sd1891, 12'sd1792}, {1'sd0, 12'sd-1673, 9'sd-210}},
{{10'sd-447, 12'sd1395, 12'sd1810}, {12'sd1649, 13'sd2770, 12'sd1854}, {11'sd606, 12'sd-1481, 9'sd-210}},
{{11'sd-973, 11'sd805, 13'sd3002}, {12'sd1337, 7'sd32, 13'sd2358}, {10'sd-310, 12'sd-1847, 11'sd-653}},
{{11'sd895, 11'sd766, 10'sd451}, {13'sd-2514, 10'sd-367, 10'sd-398}, {12'sd-1070, 11'sd696, 11'sd-774}},
{{12'sd-1556, 10'sd307, 9'sd-163}, {12'sd-2011, 12'sd-1351, 13'sd-2133}, {11'sd-927, 12'sd1307, 12'sd1288}},
{{13'sd-2383, 12'sd-1619, 13'sd-2820}, {10'sd262, 13'sd-2869, 13'sd-3016}, {4'sd6, 10'sd-369, 12'sd1556}},
{{12'sd-1755, 12'sd-1714, 13'sd-2185}, {11'sd-797, 11'sd834, 11'sd-643}, {13'sd2142, 11'sd-834, 12'sd1208}},
{{13'sd-2587, 13'sd-3882, 12'sd1608}, {13'sd-2076, 12'sd1725, 12'sd1360}, {14'sd4725, 13'sd3978, 14'sd4990}},
{{12'sd-1503, 7'sd-33, 4'sd-7}, {13'sd-2070, 12'sd-1346, 9'sd204}, {12'sd-1920, 13'sd2440, 9'sd-211}},
{{12'sd1628, 12'sd1845, 13'sd2382}, {13'sd2334, 12'sd1199, 11'sd-925}, {10'sd-270, 13'sd-2731, 12'sd1402}},
{{11'sd-744, 8'sd-115, 9'sd-191}, {11'sd932, 13'sd-2978, 12'sd-1065}, {13'sd3013, 13'sd2531, 13'sd-2777}},
{{12'sd-1615, 13'sd-3424, 9'sd-205}, {13'sd-3394, 10'sd268, 13'sd2313}, {11'sd873, 12'sd-1910, 13'sd-2202}},
{{13'sd-2927, 8'sd64, 12'sd-1200}, {13'sd-3570, 11'sd-728, 11'sd936}, {11'sd-652, 8'sd-72, 11'sd1022}},
{{13'sd3395, 13'sd3759, 13'sd2206}, {11'sd-612, 12'sd1956, 10'sd-415}, {11'sd880, 12'sd-1401, 11'sd-760}},
{{11'sd886, 12'sd-1826, 10'sd-394}, {9'sd-134, 12'sd-1614, 11'sd817}, {12'sd1216, 11'sd-558, 9'sd-198}},
{{12'sd1557, 12'sd1828, 8'sd-85}, {11'sd-968, 13'sd2283, 11'sd-637}, {13'sd-2417, 12'sd-1690, 12'sd1087}},
{{13'sd-3089, 11'sd-706, 12'sd-1356}, {12'sd1315, 10'sd-495, 13'sd-2077}, {10'sd-303, 9'sd234, 10'sd-397}},
{{11'sd-788, 12'sd1439, 12'sd-1518}, {10'sd-335, 13'sd2729, 13'sd-2602}, {11'sd851, 12'sd-1197, 12'sd-1532}},
{{12'sd1690, 13'sd2738, 11'sd582}, {13'sd-2610, 11'sd1021, 11'sd-871}, {13'sd-2393, 9'sd154, 11'sd-761}}},
{
{{12'sd-1457, 13'sd2178, 10'sd-450}, {11'sd-776, 10'sd-384, 13'sd2475}, {11'sd-771, 12'sd1386, 10'sd-434}},
{{10'sd433, 13'sd-2098, 12'sd1093}, {12'sd1493, 10'sd419, 13'sd-2540}, {11'sd547, 11'sd656, 13'sd2104}},
{{13'sd3872, 11'sd524, 11'sd806}, {11'sd-543, 12'sd-1323, 13'sd-3306}, {10'sd502, 13'sd-3228, 11'sd921}},
{{11'sd-620, 12'sd1592, 10'sd-498}, {12'sd-1664, 7'sd-50, 10'sd-262}, {11'sd-676, 9'sd157, 6'sd28}},
{{13'sd2093, 12'sd-1586, 12'sd1643}, {13'sd-2573, 12'sd1569, 13'sd2500}, {13'sd2428, 13'sd-2281, 12'sd1736}},
{{13'sd-2582, 10'sd-378, 11'sd-608}, {12'sd-1458, 10'sd410, 13'sd-2243}, {11'sd799, 12'sd-2026, 13'sd2481}},
{{13'sd2296, 11'sd-604, 13'sd-2200}, {10'sd379, 13'sd2118, 11'sd-540}, {11'sd-857, 13'sd-2328, 12'sd1906}},
{{11'sd-723, 13'sd2455, 12'sd-1514}, {10'sd408, 10'sd-315, 12'sd1512}, {12'sd1694, 13'sd2388, 11'sd638}},
{{10'sd-504, 13'sd2552, 11'sd789}, {12'sd1144, 13'sd-2180, 12'sd1121}, {13'sd-2572, 6'sd28, 13'sd-2320}},
{{13'sd2690, 12'sd-1450, 12'sd-1445}, {12'sd-1857, 6'sd25, 12'sd1698}, {10'sd-398, 10'sd-350, 12'sd1766}},
{{10'sd-489, 11'sd-596, 11'sd601}, {13'sd-2488, 13'sd-2227, 13'sd2691}, {13'sd-2910, 12'sd1404, 13'sd3762}},
{{13'sd-2485, 13'sd-2521, 13'sd-2533}, {9'sd-176, 11'sd715, 12'sd-1529}, {11'sd583, 12'sd1616, 10'sd-436}},
{{9'sd-185, 12'sd-1484, 13'sd-3129}, {12'sd-1131, 13'sd2649, 12'sd-2008}, {12'sd-1648, 13'sd2959, 11'sd943}},
{{13'sd-2831, 12'sd-1815, 12'sd1990}, {12'sd1147, 12'sd1995, 12'sd1894}, {12'sd-1843, 11'sd-854, 12'sd-1615}},
{{12'sd1879, 12'sd-2047, 11'sd674}, {10'sd-328, 12'sd-1260, 12'sd1642}, {8'sd122, 11'sd729, 10'sd-324}},
{{12'sd1560, 12'sd-1413, 12'sd-1500}, {13'sd2381, 13'sd2650, 11'sd-727}, {12'sd1735, 11'sd719, 13'sd-2681}},
{{11'sd840, 9'sd-167, 8'sd-95}, {12'sd-1806, 12'sd1850, 12'sd1312}, {13'sd3370, 11'sd-665, 13'sd2458}},
{{13'sd3880, 13'sd3333, 9'sd240}, {10'sd271, 10'sd380, 13'sd2684}, {12'sd-1062, 13'sd-3565, 13'sd-2970}},
{{11'sd-792, 12'sd-1617, 13'sd2181}, {10'sd-479, 13'sd-2294, 10'sd-323}, {10'sd331, 11'sd-577, 11'sd-1023}},
{{12'sd-1910, 11'sd-549, 13'sd2286}, {13'sd-2379, 11'sd514, 11'sd890}, {11'sd-796, 10'sd-359, 12'sd1200}},
{{12'sd1189, 13'sd2961, 12'sd-1520}, {12'sd1688, 11'sd-735, 12'sd-1607}, {12'sd1700, 13'sd-2137, 12'sd-1124}},
{{12'sd-1032, 11'sd-870, 12'sd-2012}, {11'sd-917, 5'sd13, 12'sd-1386}, {13'sd2418, 11'sd-767, 11'sd728}},
{{13'sd3031, 13'sd2833, 9'sd217}, {13'sd2471, 12'sd-1889, 10'sd-500}, {10'sd479, 12'sd1059, 12'sd-1685}},
{{11'sd-1007, 13'sd2840, 12'sd-1387}, {12'sd-1245, 13'sd2132, 12'sd-1669}, {9'sd-145, 9'sd-222, 11'sd-698}},
{{12'sd1448, 9'sd246, 10'sd348}, {13'sd2623, 13'sd2767, 13'sd-2221}, {10'sd465, 13'sd-2802, 11'sd618}},
{{12'sd-1965, 12'sd-1375, 13'sd-2499}, {12'sd-1232, 11'sd-804, 11'sd-715}, {13'sd-2266, 13'sd2654, 11'sd-749}},
{{9'sd-156, 12'sd-1349, 11'sd-896}, {13'sd-2950, 12'sd1656, 13'sd2390}, {13'sd2129, 13'sd-2889, 11'sd611}},
{{13'sd-2638, 13'sd-2461, 12'sd-1260}, {11'sd705, 11'sd-813, 12'sd-2017}, {13'sd2282, 12'sd1774, 11'sd-711}},
{{13'sd-2156, 11'sd-700, 9'sd148}, {10'sd304, 10'sd489, 13'sd-2594}, {13'sd2693, 12'sd1573, 13'sd2775}},
{{10'sd454, 13'sd-2488, 12'sd1379}, {13'sd2469, 8'sd119, 13'sd2053}, {11'sd554, 11'sd-845, 9'sd204}},
{{12'sd-1860, 9'sd244, 12'sd1549}, {11'sd-548, 12'sd-1115, 11'sd-518}, {12'sd1965, 12'sd1439, 11'sd-561}},
{{11'sd829, 11'sd-762, 13'sd2350}, {9'sd-225, 12'sd1431, 13'sd2909}, {13'sd-2424, 12'sd1321, 11'sd-633}},
{{12'sd-1275, 13'sd2264, 13'sd2465}, {12'sd-1818, 11'sd997, 12'sd-1820}, {10'sd470, 12'sd-1347, 13'sd-2393}},
{{13'sd2376, 10'sd456, 11'sd-800}, {11'sd-921, 12'sd1308, 13'sd2079}, {12'sd1400, 11'sd515, 13'sd2355}},
{{12'sd1042, 13'sd-2922, 12'sd-1887}, {11'sd-788, 11'sd-1010, 12'sd1173}, {11'sd925, 13'sd-2290, 8'sd-103}},
{{12'sd-1536, 13'sd-2457, 10'sd-462}, {9'sd-240, 11'sd770, 13'sd-2771}, {10'sd-444, 12'sd1080, 13'sd-2395}},
{{12'sd-1480, 11'sd793, 11'sd-756}, {10'sd-286, 7'sd62, 11'sd642}, {8'sd-114, 12'sd-1363, 12'sd-1981}},
{{12'sd1493, 13'sd-2126, 10'sd-419}, {8'sd-86, 7'sd-58, 11'sd-808}, {11'sd-814, 13'sd3007, 13'sd2282}},
{{9'sd162, 13'sd-2372, 12'sd1354}, {13'sd2587, 12'sd1698, 13'sd-2153}, {13'sd3721, 12'sd1176, 13'sd2071}},
{{13'sd-2638, 12'sd-1230, 12'sd-1207}, {12'sd1042, 12'sd1612, 12'sd-1887}, {13'sd2845, 10'sd439, 12'sd-1479}},
{{10'sd-343, 12'sd1845, 11'sd640}, {11'sd721, 13'sd-2115, 10'sd456}, {13'sd-2513, 13'sd-2217, 11'sd991}},
{{11'sd-785, 11'sd772, 11'sd-785}, {13'sd-2067, 12'sd-1230, 10'sd316}, {10'sd418, 11'sd-908, 10'sd-308}},
{{9'sd-175, 12'sd-1654, 10'sd-413}, {12'sd1775, 12'sd-1140, 11'sd954}, {11'sd-796, 13'sd2115, 10'sd321}},
{{11'sd751, 10'sd-360, 9'sd-225}, {13'sd-3480, 13'sd-2232, 12'sd-1273}, {12'sd-1715, 9'sd170, 12'sd-1790}},
{{10'sd443, 13'sd2606, 13'sd-2608}, {13'sd-2707, 9'sd212, 12'sd-1919}, {10'sd-471, 8'sd72, 12'sd-1700}},
{{12'sd1074, 11'sd-584, 11'sd800}, {11'sd-630, 11'sd676, 9'sd246}, {9'sd197, 11'sd-519, 11'sd-761}},
{{13'sd2485, 12'sd1379, 11'sd1003}, {13'sd3380, 10'sd-267, 13'sd-2671}, {11'sd790, 12'sd1354, 11'sd929}},
{{12'sd1689, 13'sd2390, 13'sd-2682}, {12'sd-1692, 11'sd-534, 7'sd-63}, {11'sd772, 10'sd-498, 11'sd660}},
{{13'sd-2657, 12'sd1853, 11'sd-1009}, {9'sd170, 11'sd-661, 11'sd973}, {8'sd123, 10'sd-424, 13'sd2510}},
{{11'sd-978, 12'sd1102, 13'sd2049}, {11'sd1019, 11'sd-907, 11'sd945}, {12'sd1683, 12'sd1276, 12'sd-1855}},
{{13'sd-2513, 11'sd918, 12'sd1598}, {11'sd-745, 13'sd2098, 13'sd-2437}, {11'sd-780, 12'sd1704, 12'sd1426}},
{{13'sd-2679, 11'sd-711, 12'sd-1969}, {12'sd-1383, 12'sd2041, 13'sd2072}, {13'sd-2212, 10'sd-346, 11'sd-626}},
{{12'sd1270, 10'sd428, 13'sd2523}, {12'sd-1195, 9'sd-160, 13'sd2121}, {13'sd-2505, 13'sd-2918, 6'sd-22}},
{{12'sd1802, 13'sd2896, 11'sd594}, {13'sd3046, 12'sd1656, 12'sd1275}, {9'sd143, 9'sd243, 12'sd-1916}},
{{13'sd2963, 11'sd1001, 8'sd-120}, {13'sd2956, 12'sd1065, 11'sd-770}, {13'sd2948, 12'sd1237, 13'sd2392}},
{{13'sd2264, 13'sd-2411, 12'sd1342}, {12'sd-1335, 7'sd-50, 10'sd-262}, {12'sd1636, 8'sd-94, 13'sd-2205}},
{{12'sd1421, 13'sd2212, 12'sd-1056}, {11'sd688, 11'sd608, 12'sd1999}, {12'sd1443, 13'sd2564, 12'sd-1195}},
{{12'sd-1225, 2'sd-1, 13'sd2841}, {12'sd-1818, 12'sd-1562, 11'sd-818}, {11'sd-534, 8'sd-115, 11'sd997}},
{{12'sd1231, 13'sd3074, 11'sd-835}, {12'sd-1231, 13'sd-2529, 12'sd1784}, {12'sd-1358, 13'sd-3474, 9'sd-155}},
{{13'sd-2914, 12'sd-1521, 12'sd1872}, {12'sd1827, 13'sd-2312, 10'sd410}, {11'sd767, 12'sd1505, 12'sd-1321}},
{{12'sd1330, 13'sd2637, 11'sd-959}, {10'sd308, 11'sd-572, 13'sd-2186}, {11'sd-783, 11'sd743, 13'sd-2159}},
{{12'sd-1042, 13'sd-2989, 11'sd829}, {8'sd110, 11'sd-987, 13'sd2491}, {12'sd-1174, 12'sd-1365, 13'sd-2137}},
{{12'sd-1900, 12'sd1957, 13'sd-2663}, {13'sd-2423, 12'sd1374, 12'sd-1595}, {13'sd-2402, 13'sd2807, 11'sd995}},
{{12'sd-1313, 13'sd2088, 11'sd704}, {13'sd2643, 13'sd2535, 11'sd-613}, {11'sd756, 12'sd1672, 11'sd-769}}},
{
{{14'sd4277, 10'sd369, 13'sd2633}, {11'sd-725, 11'sd882, 12'sd-1584}, {10'sd-328, 9'sd185, 12'sd-1847}},
{{13'sd2729, 10'sd-474, 9'sd-184}, {9'sd201, 12'sd1822, 13'sd-2440}, {12'sd1463, 12'sd-1633, 13'sd-2551}},
{{13'sd3881, 13'sd3668, 12'sd-1899}, {10'sd426, 14'sd4441, 9'sd-232}, {6'sd21, 11'sd637, 11'sd-615}},
{{8'sd89, 12'sd-2000, 12'sd1226}, {12'sd-1583, 11'sd-577, 9'sd167}, {12'sd1606, 12'sd-1198, 13'sd2097}},
{{14'sd4711, 13'sd-2792, 12'sd-1189}, {11'sd-981, 12'sd-1921, 13'sd2452}, {10'sd356, 9'sd177, 12'sd-1808}},
{{12'sd-1104, 13'sd-2508, 10'sd-332}, {12'sd-1418, 12'sd-1175, 13'sd-2208}, {10'sd-400, 13'sd-2048, 11'sd-745}},
{{10'sd266, 13'sd2078, 13'sd2286}, {12'sd1074, 13'sd-2391, 13'sd2220}, {12'sd1283, 11'sd541, 12'sd1048}},
{{12'sd-1649, 11'sd-706, 11'sd699}, {12'sd-1162, 12'sd-1636, 13'sd-2184}, {11'sd-681, 12'sd1680, 10'sd-442}},
{{12'sd-1778, 13'sd-3166, 11'sd-843}, {13'sd-3140, 10'sd-262, 12'sd1740}, {11'sd681, 13'sd-2100, 10'sd280}},
{{11'sd-620, 12'sd-1575, 12'sd1762}, {14'sd4171, 12'sd-1702, 11'sd644}, {13'sd3278, 11'sd944, 13'sd2739}},
{{13'sd-3804, 14'sd-4105, 11'sd-598}, {11'sd977, 13'sd-3410, 10'sd-423}, {12'sd-1479, 11'sd-536, 12'sd-1052}},
{{10'sd272, 10'sd345, 12'sd1387}, {12'sd-1505, 13'sd-2847, 13'sd2404}, {12'sd-1312, 13'sd2475, 12'sd1304}},
{{13'sd-3149, 13'sd3095, 13'sd-3105}, {13'sd-3821, 11'sd1017, 13'sd-2763}, {11'sd-683, 12'sd-1156, 13'sd2686}},
{{12'sd-1263, 13'sd-2346, 11'sd824}, {11'sd516, 12'sd-1037, 13'sd-2574}, {13'sd2412, 12'sd1971, 12'sd1170}},
{{11'sd-537, 9'sd-209, 13'sd2806}, {9'sd214, 13'sd-2214, 10'sd-279}, {12'sd-1151, 12'sd-1655, 11'sd-559}},
{{9'sd226, 12'sd1989, 12'sd1385}, {13'sd3181, 12'sd-1679, 13'sd-2108}, {13'sd3961, 12'sd-1526, 13'sd-2071}},
{{11'sd-958, 13'sd3702, 12'sd1203}, {13'sd-2055, 12'sd-1959, 11'sd-835}, {13'sd-2295, 11'sd551, 13'sd2181}},
{{14'sd6897, 14'sd4537, 12'sd1709}, {14'sd4938, 11'sd-598, 12'sd-1033}, {13'sd2387, 12'sd1494, 13'sd-3592}},
{{11'sd667, 13'sd2305, 13'sd2837}, {12'sd1752, 13'sd-2186, 12'sd-1112}, {12'sd-1538, 12'sd-1516, 12'sd-1261}},
{{13'sd-3645, 11'sd-1018, 13'sd2370}, {12'sd1188, 13'sd-2600, 11'sd-912}, {11'sd-874, 13'sd-2318, 12'sd-1062}},
{{13'sd2503, 11'sd-644, 12'sd1107}, {10'sd442, 12'sd-1538, 12'sd-1084}, {10'sd274, 12'sd1195, 12'sd-1885}},
{{13'sd3885, 12'sd1876, 12'sd1942}, {12'sd1885, 13'sd2105, 11'sd-576}, {12'sd-1712, 13'sd-2707, 11'sd-636}},
{{12'sd-1207, 10'sd-386, 9'sd-239}, {12'sd1574, 11'sd594, 12'sd-1624}, {13'sd2561, 12'sd-1845, 13'sd2730}},
{{12'sd1703, 13'sd2557, 12'sd1693}, {10'sd256, 10'sd-497, 13'sd2526}, {13'sd-2449, 13'sd2338, 13'sd2829}},
{{12'sd-1487, 11'sd-627, 12'sd-1890}, {11'sd929, 12'sd1335, 13'sd-2069}, {13'sd2589, 13'sd3543, 12'sd1752}},
{{12'sd1179, 8'sd105, 11'sd523}, {12'sd1094, 11'sd1014, 12'sd-1681}, {10'sd378, 11'sd-522, 13'sd-2095}},
{{12'sd-1250, 12'sd-1762, 12'sd1558}, {12'sd1471, 12'sd1042, 11'sd-832}, {13'sd-2448, 10'sd344, 13'sd2633}},
{{12'sd-1551, 11'sd-876, 12'sd1643}, {12'sd-1778, 13'sd-2588, 11'sd658}, {13'sd2433, 12'sd-1186, 11'sd628}},
{{9'sd-205, 9'sd-147, 10'sd256}, {13'sd-2962, 12'sd1412, 13'sd2634}, {13'sd-2263, 13'sd-3119, 13'sd-2782}},
{{9'sd191, 13'sd2216, 10'sd509}, {12'sd-1045, 10'sd492, 12'sd-1111}, {11'sd879, 10'sd-482, 10'sd480}},
{{13'sd-2671, 12'sd-1798, 11'sd704}, {10'sd-440, 12'sd1960, 12'sd1640}, {13'sd-3745, 11'sd-870, 11'sd-900}},
{{12'sd-1528, 11'sd-767, 12'sd1107}, {11'sd-981, 9'sd-140, 10'sd410}, {13'sd3202, 13'sd-2586, 12'sd-1300}},
{{10'sd307, 12'sd-1640, 12'sd1835}, {11'sd973, 11'sd-971, 10'sd480}, {13'sd-2091, 13'sd-2072, 12'sd-1818}},
{{12'sd-1568, 12'sd1652, 13'sd2772}, {11'sd-669, 11'sd-690, 10'sd-361}, {10'sd-406, 11'sd-1016, 11'sd-691}},
{{12'sd-1445, 13'sd2161, 11'sd-863}, {12'sd-1899, 10'sd-350, 12'sd2032}, {12'sd-1291, 12'sd-1420, 12'sd-1749}},
{{12'sd-2045, 8'sd104, 13'sd-2772}, {13'sd2396, 12'sd1884, 10'sd396}, {12'sd1233, 11'sd559, 9'sd-244}},
{{11'sd-522, 13'sd2964, 12'sd-1212}, {13'sd-2980, 12'sd1614, 13'sd-2974}, {10'sd461, 12'sd1600, 12'sd1094}},
{{13'sd3984, 12'sd1831, 13'sd-2657}, {14'sd5937, 13'sd-2523, 13'sd-2221}, {14'sd5263, 12'sd-1433, 13'sd-3600}},
{{12'sd-1775, 13'sd-2327, 13'sd-2477}, {13'sd3526, 10'sd360, 11'sd-775}, {14'sd4109, 11'sd584, 5'sd-13}},
{{8'sd-80, 13'sd-2511, 10'sd317}, {6'sd-16, 13'sd-3037, 10'sd-317}, {13'sd2214, 12'sd-1594, 13'sd-3460}},
{{12'sd1468, 13'sd-2442, 12'sd-1375}, {13'sd2596, 11'sd956, 13'sd-2091}, {11'sd652, 11'sd756, 13'sd-2432}},
{{11'sd920, 12'sd1559, 10'sd466}, {12'sd-1186, 12'sd-1736, 13'sd-2579}, {10'sd-332, 13'sd2540, 13'sd2725}},
{{13'sd-2588, 11'sd-530, 12'sd1127}, {12'sd2009, 11'sd-626, 13'sd-2135}, {11'sd-529, 13'sd-2318, 12'sd-1052}},
{{13'sd-2086, 11'sd-996, 10'sd285}, {14'sd-5091, 12'sd2007, 12'sd-1353}, {13'sd-3472, 13'sd-2380, 14'sd4389}},
{{12'sd-1370, 9'sd-172, 13'sd3163}, {13'sd2178, 12'sd1121, 12'sd1736}, {13'sd-3075, 13'sd2108, 12'sd1374}},
{{13'sd3023, 8'sd-100, 12'sd1837}, {12'sd1091, 9'sd167, 12'sd-1340}, {13'sd2452, 13'sd2231, 12'sd-2026}},
{{14'sd4579, 12'sd-1388, 12'sd-1399}, {11'sd941, 3'sd2, 13'sd-2979}, {12'sd-1263, 13'sd2436, 11'sd-711}},
{{11'sd787, 12'sd1797, 13'sd2374}, {12'sd1739, 10'sd341, 13'sd2765}, {12'sd-1237, 13'sd-2418, 8'sd-78}},
{{8'sd67, 13'sd-2567, 5'sd13}, {8'sd83, 12'sd-1048, 12'sd1218}, {12'sd-1542, 12'sd1190, 13'sd2268}},
{{12'sd-1722, 13'sd2454, 13'sd2366}, {12'sd1568, 11'sd589, 11'sd-630}, {12'sd-1681, 9'sd155, 13'sd-2386}},
{{10'sd-367, 13'sd3098, 12'sd-1734}, {12'sd-1837, 9'sd230, 12'sd1161}, {9'sd-232, 12'sd-1570, 13'sd-2557}},
{{13'sd2156, 12'sd-1140, 12'sd1493}, {9'sd184, 12'sd1875, 13'sd2531}, {12'sd1581, 11'sd-754, 10'sd-460}},
{{13'sd3926, 12'sd-1248, 11'sd604}, {12'sd1885, 9'sd-147, 12'sd-1308}, {12'sd1633, 13'sd-2587, 11'sd-825}},
{{9'sd-246, 11'sd890, 12'sd1899}, {12'sd-1505, 12'sd1641, 12'sd-1966}, {12'sd1297, 12'sd1389, 12'sd-1522}},
{{12'sd-1793, 13'sd2605, 12'sd1410}, {11'sd-822, 12'sd-1825, 9'sd185}, {12'sd1900, 13'sd2417, 10'sd-280}},
{{13'sd-2581, 9'sd180, 12'sd2041}, {9'sd231, 10'sd325, 12'sd-1288}, {12'sd1967, 11'sd-915, 12'sd-1829}},
{{13'sd-2681, 12'sd1674, 10'sd-323}, {13'sd-2609, 12'sd-1486, 6'sd24}, {12'sd1131, 12'sd-1639, 7'sd47}},
{{11'sd-566, 12'sd-1362, 11'sd613}, {11'sd636, 13'sd-3807, 13'sd3137}, {12'sd1506, 11'sd892, 11'sd-737}},
{{12'sd-1123, 13'sd-3460, 13'sd2366}, {12'sd-1692, 13'sd2210, 13'sd3409}, {12'sd2011, 11'sd562, 8'sd-111}},
{{13'sd2951, 13'sd2290, 12'sd-2008}, {11'sd633, 12'sd1372, 12'sd-1965}, {13'sd2890, 13'sd-2474, 11'sd776}},
{{11'sd-620, 9'sd199, 13'sd-3236}, {10'sd498, 12'sd1402, 12'sd1486}, {13'sd3522, 12'sd-1285, 10'sd-406}},
{{10'sd-507, 12'sd1392, 13'sd2322}, {11'sd832, 13'sd-2406, 12'sd-1806}, {12'sd1519, 13'sd2718, 11'sd-601}},
{{12'sd-1444, 13'sd-2515, 12'sd1791}, {12'sd-1778, 10'sd-314, 12'sd-1578}, {13'sd-2397, 13'sd-2386, 12'sd1803}},
{{13'sd3069, 13'sd-2166, 11'sd-850}, {11'sd-921, 13'sd-2466, 12'sd1840}, {11'sd600, 13'sd-2558, 11'sd753}}},
{
{{11'sd-1018, 12'sd-1890, 12'sd-1107}, {11'sd-592, 9'sd252, 13'sd3626}, {12'sd-1335, 10'sd-423, 12'sd1744}},
{{11'sd-660, 12'sd1682, 13'sd-2470}, {12'sd1389, 12'sd1556, 13'sd-3232}, {13'sd-3103, 12'sd-1939, 8'sd-105}},
{{9'sd222, 12'sd1080, 13'sd-2524}, {12'sd1556, 13'sd2805, 11'sd916}, {12'sd-1910, 12'sd-2030, 12'sd1405}},
{{12'sd1525, 12'sd1975, 11'sd743}, {13'sd2888, 10'sd-363, 12'sd-1224}, {12'sd1971, 11'sd-982, 12'sd1613}},
{{13'sd-2993, 12'sd1867, 10'sd473}, {13'sd-2195, 11'sd-643, 12'sd1284}, {12'sd-1306, 11'sd-777, 10'sd350}},
{{11'sd-581, 12'sd1223, 13'sd2751}, {8'sd-93, 13'sd-2767, 8'sd70}, {12'sd-1326, 12'sd1589, 12'sd1037}},
{{10'sd-387, 12'sd-1083, 12'sd-1995}, {12'sd1894, 12'sd-1907, 12'sd2024}, {12'sd1819, 12'sd1235, 13'sd3237}},
{{10'sd-458, 11'sd700, 13'sd-3122}, {12'sd-1081, 12'sd1286, 10'sd-381}, {13'sd-2314, 9'sd-236, 10'sd-503}},
{{13'sd-2543, 13'sd-2231, 13'sd-2387}, {13'sd-3213, 11'sd968, 13'sd-2788}, {11'sd-647, 13'sd-2200, 13'sd-3593}},
{{11'sd889, 10'sd-408, 13'sd-2230}, {12'sd1630, 12'sd-1528, 12'sd-1553}, {13'sd-2235, 10'sd-316, 11'sd930}},
{{11'sd934, 12'sd1511, 14'sd4669}, {13'sd2186, 9'sd218, 11'sd946}, {12'sd-1778, 13'sd-2273, 12'sd1694}},
{{13'sd2996, 12'sd1868, 12'sd1377}, {12'sd-1031, 10'sd495, 7'sd34}, {13'sd-3177, 10'sd390, 13'sd-2756}},
{{11'sd-853, 7'sd-32, 11'sd-852}, {13'sd2451, 12'sd1077, 10'sd451}, {12'sd-1231, 11'sd-609, 11'sd-641}},
{{12'sd-1823, 12'sd1092, 13'sd-2850}, {13'sd2804, 10'sd456, 12'sd-1027}, {11'sd-823, 9'sd-225, 13'sd-3196}},
{{11'sd-959, 11'sd1004, 12'sd-1783}, {12'sd1192, 13'sd2170, 9'sd146}, {12'sd-1621, 13'sd2192, 12'sd-1974}},
{{7'sd-51, 10'sd502, 10'sd285}, {13'sd-2920, 12'sd1622, 12'sd-1183}, {9'sd-171, 13'sd2277, 11'sd748}},
{{14'sd4981, 10'sd-347, 10'sd-273}, {11'sd-991, 8'sd-117, 13'sd-2394}, {11'sd593, 13'sd3387, 10'sd-273}},
{{14'sd-4157, 14'sd-5769, 14'sd-5587}, {12'sd1125, 12'sd-1192, 11'sd924}, {9'sd224, 13'sd2944, 13'sd2602}},
{{6'sd-21, 12'sd-1708, 13'sd-2768}, {13'sd2592, 13'sd-2193, 9'sd220}, {12'sd-1240, 12'sd-1264, 12'sd-1786}},
{{9'sd147, 8'sd113, 14'sd-5013}, {12'sd1778, 11'sd973, 12'sd-1594}, {13'sd2727, 11'sd-535, 13'sd-2166}},
{{12'sd-1399, 13'sd-2295, 12'sd1341}, {12'sd1333, 13'sd-2452, 10'sd-493}, {12'sd1438, 13'sd-2210, 12'sd-1430}},
{{13'sd-3360, 13'sd-3704, 11'sd1011}, {12'sd-1993, 12'sd1186, 8'sd92}, {13'sd-2271, 9'sd-231, 12'sd-1278}},
{{10'sd370, 13'sd-2893, 13'sd2874}, {13'sd-2141, 13'sd2130, 11'sd953}, {12'sd-1924, 10'sd421, 12'sd1345}},
{{12'sd1153, 9'sd169, 11'sd-1014}, {13'sd-2434, 12'sd1033, 13'sd-2751}, {7'sd42, 13'sd-2315, 5'sd11}},
{{13'sd2844, 14'sd4735, 11'sd993}, {12'sd1037, 13'sd3848, 13'sd3181}, {12'sd1572, 11'sd-572, 13'sd2682}},
{{10'sd321, 11'sd-987, 13'sd-2628}, {9'sd-134, 12'sd1450, 13'sd2257}, {12'sd-1720, 11'sd1022, 12'sd1736}},
{{12'sd1841, 12'sd1982, 8'sd100}, {11'sd546, 11'sd-812, 12'sd1553}, {10'sd-497, 12'sd1325, 9'sd134}},
{{13'sd2416, 12'sd1822, 11'sd659}, {11'sd953, 13'sd2592, 11'sd565}, {9'sd-229, 12'sd-1773, 12'sd1495}},
{{11'sd935, 13'sd-3660, 12'sd-1096}, {13'sd2556, 13'sd-2208, 12'sd-1367}, {11'sd739, 12'sd2005, 13'sd2330}},
{{13'sd-2126, 12'sd-1469, 9'sd142}, {13'sd-2256, 7'sd63, 11'sd-615}, {13'sd2370, 10'sd-428, 9'sd-182}},
{{11'sd632, 11'sd-1018, 12'sd1295}, {12'sd-1133, 11'sd755, 12'sd1584}, {11'sd974, 12'sd1215, 10'sd468}},
{{13'sd-2367, 12'sd-1858, 13'sd-4012}, {13'sd2685, 13'sd2355, 13'sd-2272}, {12'sd-1571, 11'sd-982, 10'sd497}},
{{13'sd-2738, 12'sd-1113, 13'sd-3258}, {13'sd2577, 12'sd1131, 13'sd2772}, {8'sd103, 13'sd2837, 13'sd3448}},
{{11'sd733, 11'sd541, 11'sd-999}, {12'sd-1959, 12'sd-1090, 12'sd1784}, {12'sd-1987, 13'sd-2427, 13'sd3186}},
{{12'sd1446, 11'sd903, 8'sd71}, {12'sd-1085, 11'sd-902, 13'sd-2915}, {10'sd472, 12'sd1656, 12'sd1744}},
{{13'sd2430, 11'sd756, 10'sd437}, {12'sd-1823, 12'sd-1680, 9'sd-138}, {10'sd481, 10'sd-498, 13'sd-3354}},
{{12'sd-1900, 11'sd966, 13'sd-2923}, {13'sd-3104, 12'sd1422, 13'sd-3225}, {12'sd-1578, 12'sd-2001, 12'sd1659}},
{{9'sd-178, 10'sd389, 12'sd-1847}, {13'sd-2860, 9'sd244, 11'sd-678}, {13'sd-4018, 13'sd2606, 11'sd813}},
{{13'sd3624, 11'sd799, 12'sd-1586}, {13'sd2085, 11'sd578, 11'sd-1018}, {13'sd2380, 11'sd-1023, 9'sd-217}},
{{11'sd613, 11'sd1014, 10'sd266}, {12'sd-1094, 12'sd1444, 12'sd1474}, {13'sd-3070, 13'sd2232, 12'sd2004}},
{{12'sd-1732, 8'sd100, 12'sd1237}, {11'sd895, 11'sd765, 10'sd480}, {13'sd2394, 11'sd-745, 12'sd1245}},
{{11'sd-732, 13'sd2929, 12'sd-1505}, {13'sd-2582, 12'sd1935, 9'sd-212}, {11'sd932, 12'sd-1346, 13'sd-2875}},
{{12'sd1478, 12'sd1312, 10'sd-500}, {13'sd-2091, 11'sd-694, 12'sd-1904}, {12'sd-2011, 11'sd-978, 13'sd-3481}},
{{11'sd-738, 12'sd-1330, 12'sd1442}, {10'sd430, 10'sd424, 10'sd-464}, {12'sd-1419, 11'sd837, 11'sd-962}},
{{13'sd-3520, 11'sd866, 6'sd-23}, {11'sd-557, 13'sd-2618, 12'sd-1093}, {11'sd-723, 13'sd-2417, 10'sd-496}},
{{14'sd-4944, 13'sd-3590, 10'sd257}, {13'sd-2461, 10'sd-499, 12'sd1127}, {13'sd-2989, 11'sd-786, 12'sd1582}},
{{13'sd2235, 13'sd2372, 13'sd-2544}, {11'sd-743, 11'sd-1016, 13'sd2782}, {13'sd2853, 11'sd-538, 14'sd4746}},
{{13'sd-2730, 11'sd808, 12'sd-1452}, {12'sd1612, 12'sd-2043, 12'sd-1275}, {9'sd255, 12'sd-1967, 13'sd-2573}},
{{12'sd-1350, 12'sd1062, 13'sd-3302}, {12'sd1903, 7'sd37, 13'sd2144}, {13'sd2712, 10'sd-260, 13'sd-2282}},
{{11'sd-1001, 9'sd241, 13'sd3445}, {11'sd-749, 12'sd-1199, 12'sd1388}, {13'sd-2093, 13'sd3253, 11'sd704}},
{{6'sd18, 10'sd-469, 10'sd-341}, {10'sd-401, 11'sd655, 13'sd-2073}, {11'sd885, 12'sd1854, 9'sd186}},
{{12'sd1087, 13'sd2550, 12'sd-1138}, {12'sd-1511, 12'sd-1728, 12'sd-1425}, {11'sd675, 5'sd-10, 13'sd2121}},
{{11'sd873, 12'sd-1290, 13'sd2310}, {8'sd-94, 9'sd136, 7'sd-50}, {11'sd-574, 11'sd-817, 12'sd1981}},
{{10'sd256, 13'sd2361, 11'sd-806}, {8'sd-106, 13'sd-2444, 13'sd3041}, {12'sd-1532, 13'sd2925, 12'sd-1579}},
{{12'sd-1587, 13'sd2360, 10'sd296}, {12'sd-1502, 12'sd-1293, 8'sd-113}, {13'sd2701, 12'sd-1727, 13'sd3404}},
{{13'sd-3211, 12'sd-1422, 13'sd2782}, {12'sd-1965, 10'sd-375, 9'sd168}, {12'sd1288, 12'sd-1862, 10'sd266}},
{{12'sd1808, 12'sd1143, 13'sd2480}, {7'sd-52, 13'sd2247, 13'sd2627}, {13'sd2121, 12'sd1911, 12'sd-1453}},
{{11'sd-898, 10'sd-437, 11'sd-1009}, {12'sd-1445, 6'sd25, 11'sd-854}, {12'sd-1877, 12'sd1568, 11'sd775}},
{{12'sd-1433, 7'sd34, 13'sd-3617}, {13'sd-2070, 10'sd-444, 13'sd-2281}, {12'sd2010, 10'sd-420, 10'sd-263}},
{{13'sd2515, 11'sd-513, 13'sd-2718}, {12'sd-1289, 12'sd-2011, 12'sd-1854}, {9'sd-136, 12'sd-1173, 12'sd-1732}},
{{12'sd-1813, 13'sd2685, 11'sd530}, {12'sd-1920, 12'sd-1795, 7'sd-56}, {6'sd-26, 12'sd1157, 11'sd-796}},
{{13'sd3991, 12'sd1284, 12'sd-1170}, {13'sd-2137, 13'sd2815, 10'sd382}, {12'sd-1506, 13'sd-2380, 12'sd-1859}},
{{13'sd-3056, 12'sd1187, 11'sd1012}, {10'sd444, 13'sd-2800, 10'sd271}, {10'sd475, 5'sd11, 12'sd1036}},
{{13'sd2358, 13'sd2577, 13'sd-2844}, {12'sd-1632, 12'sd-1365, 12'sd-1352}, {11'sd980, 12'sd-1760, 13'sd2676}}},
{
{{11'sd731, 11'sd-532, 13'sd-2155}, {11'sd-916, 11'sd769, 12'sd-1262}, {12'sd2018, 12'sd1729, 13'sd-3230}},
{{11'sd800, 12'sd-1497, 12'sd-1975}, {10'sd-386, 13'sd-2532, 13'sd2408}, {12'sd-1943, 13'sd2242, 13'sd-2357}},
{{12'sd-1517, 12'sd1658, 10'sd307}, {13'sd-3285, 13'sd-2503, 9'sd-212}, {12'sd-1583, 12'sd-1045, 13'sd3218}},
{{12'sd1881, 12'sd-1990, 11'sd728}, {5'sd15, 12'sd-1186, 13'sd2721}, {11'sd931, 12'sd1937, 9'sd128}},
{{10'sd368, 13'sd2507, 11'sd-759}, {12'sd1403, 13'sd2679, 6'sd31}, {12'sd-1427, 10'sd360, 10'sd329}},
{{11'sd-608, 10'sd323, 9'sd222}, {11'sd-685, 10'sd-285, 12'sd-1372}, {8'sd-109, 11'sd549, 11'sd951}},
{{11'sd703, 13'sd-2130, 12'sd1922}, {10'sd341, 11'sd1013, 13'sd-2067}, {10'sd-377, 11'sd849, 11'sd-541}},
{{9'sd-234, 13'sd2299, 11'sd674}, {12'sd-1493, 12'sd-1421, 11'sd-694}, {13'sd-2888, 10'sd470, 12'sd1598}},
{{10'sd-335, 11'sd936, 12'sd1572}, {12'sd1128, 11'sd-804, 12'sd1175}, {10'sd490, 11'sd-819, 12'sd-1722}},
{{10'sd-447, 13'sd-2894, 11'sd-737}, {13'sd-2331, 13'sd-2683, 12'sd-1903}, {13'sd2103, 13'sd2578, 12'sd1340}},
{{13'sd3241, 10'sd-423, 12'sd-1972}, {13'sd2102, 12'sd-2016, 13'sd-3308}, {11'sd-872, 13'sd-2272, 11'sd-997}},
{{10'sd-387, 9'sd-141, 11'sd-671}, {10'sd506, 11'sd829, 13'sd2425}, {12'sd1505, 11'sd-725, 10'sd-486}},
{{13'sd2212, 8'sd73, 13'sd-2104}, {12'sd-1044, 13'sd-2257, 10'sd321}, {11'sd567, 12'sd1597, 11'sd889}},
{{11'sd632, 12'sd1134, 13'sd-2191}, {13'sd2196, 12'sd-1232, 13'sd2426}, {12'sd2003, 12'sd1764, 13'sd-2545}},
{{13'sd2512, 13'sd-2321, 10'sd-389}, {11'sd-889, 12'sd1527, 12'sd-1514}, {9'sd136, 9'sd-205, 12'sd1761}},
{{9'sd170, 10'sd429, 12'sd1921}, {11'sd910, 12'sd1163, 13'sd2613}, {13'sd-2328, 10'sd353, 12'sd1470}},
{{12'sd1948, 13'sd2468, 13'sd2262}, {12'sd1942, 12'sd1787, 11'sd665}, {12'sd1668, 11'sd583, 12'sd1141}},
{{14'sd-5801, 13'sd-3147, 5'sd9}, {9'sd-135, 13'sd-2825, 11'sd854}, {11'sd-812, 13'sd3462, 14'sd4182}},
{{10'sd-295, 13'sd2748, 12'sd-1030}, {12'sd-1264, 13'sd2183, 13'sd2543}, {12'sd1383, 4'sd5, 12'sd1794}},
{{11'sd-595, 13'sd-2334, 9'sd-177}, {12'sd-1138, 13'sd2112, 11'sd671}, {13'sd2461, 12'sd-1789, 11'sd561}},
{{11'sd-619, 13'sd-2506, 12'sd1082}, {11'sd-717, 7'sd-43, 11'sd-820}, {12'sd-1451, 12'sd-1658, 13'sd-2354}},
{{11'sd829, 13'sd2117, 12'sd2000}, {12'sd1527, 12'sd1504, 13'sd2357}, {13'sd-2374, 11'sd-711, 12'sd1901}},
{{11'sd-657, 12'sd-1467, 12'sd1563}, {12'sd-1625, 12'sd-1832, 12'sd-1940}, {12'sd-1519, 11'sd549, 12'sd-1076}},
{{12'sd-1668, 13'sd-2964, 12'sd-1469}, {11'sd830, 12'sd-1431, 12'sd1244}, {11'sd-931, 11'sd-757, 12'sd-1449}},
{{13'sd-2621, 13'sd2362, 12'sd-1122}, {6'sd30, 13'sd-2797, 7'sd-40}, {13'sd-3221, 13'sd2058, 13'sd2683}},
{{11'sd-692, 8'sd-108, 12'sd-1411}, {12'sd2047, 12'sd-1548, 11'sd987}, {13'sd-2230, 12'sd-1841, 11'sd-978}},
{{12'sd-1870, 10'sd301, 10'sd-428}, {12'sd1923, 10'sd-488, 12'sd1100}, {11'sd1014, 12'sd1345, 11'sd-688}},
{{7'sd45, 11'sd-523, 12'sd1641}, {13'sd-2597, 12'sd1505, 12'sd-1878}, {12'sd1340, 12'sd-1035, 9'sd-251}},
{{13'sd2475, 12'sd-1901, 13'sd-2769}, {12'sd1775, 13'sd-2287, 13'sd2447}, {13'sd2375, 12'sd1884, 10'sd273}},
{{12'sd1675, 11'sd873, 12'sd-1596}, {8'sd88, 11'sd746, 12'sd-1583}, {11'sd760, 12'sd1522, 13'sd2213}},
{{11'sd516, 11'sd-771, 11'sd611}, {12'sd-1867, 12'sd1627, 11'sd-688}, {11'sd-859, 11'sd731, 13'sd2456}},
{{11'sd784, 12'sd-1707, 13'sd2228}, {12'sd1484, 10'sd-314, 13'sd2088}, {13'sd-2622, 12'sd1644, 12'sd-1798}},
{{12'sd-1268, 10'sd324, 11'sd908}, {9'sd-149, 13'sd-2478, 11'sd-675}, {13'sd2435, 12'sd-1903, 12'sd2032}},
{{12'sd-1221, 7'sd38, 11'sd969}, {12'sd1375, 11'sd865, 12'sd-1798}, {12'sd-1233, 11'sd622, 12'sd-1229}},
{{10'sd-291, 12'sd1349, 12'sd2019}, {11'sd783, 12'sd1904, 12'sd-1504}, {11'sd1015, 12'sd1101, 12'sd-1536}},
{{10'sd297, 13'sd2937, 13'sd2404}, {4'sd4, 10'sd-397, 12'sd1411}, {11'sd744, 13'sd2864, 12'sd-1929}},
{{12'sd-1253, 13'sd-2804, 12'sd1089}, {12'sd-1264, 12'sd-1357, 10'sd-424}, {13'sd3216, 11'sd788, 11'sd900}},
{{12'sd1401, 12'sd1589, 12'sd-2011}, {12'sd1096, 13'sd2266, 13'sd-2474}, {13'sd-2465, 11'sd-842, 10'sd-418}},
{{11'sd571, 11'sd-524, 12'sd1323}, {11'sd-606, 12'sd1085, 12'sd-1391}, {13'sd2140, 12'sd-1379, 12'sd-1764}},
{{12'sd1259, 13'sd2757, 12'sd-1575}, {13'sd-2073, 11'sd681, 12'sd-1425}, {12'sd-1746, 11'sd526, 12'sd-1027}},
{{12'sd-1253, 11'sd907, 13'sd-2218}, {12'sd-1919, 10'sd333, 11'sd680}, {13'sd-2312, 12'sd-1092, 11'sd-613}},
{{12'sd1749, 12'sd1456, 13'sd-2180}, {12'sd-1934, 11'sd-679, 11'sd1000}, {12'sd1785, 13'sd2170, 12'sd-1241}},
{{13'sd2155, 6'sd19, 11'sd-747}, {12'sd1631, 10'sd-281, 12'sd-1564}, {12'sd1349, 13'sd2307, 12'sd1146}},
{{10'sd285, 11'sd723, 12'sd1793}, {13'sd2777, 10'sd-262, 10'sd511}, {11'sd-642, 6'sd-24, 11'sd-815}},
{{12'sd-1452, 9'sd-212, 12'sd2039}, {9'sd219, 12'sd-1589, 12'sd-1845}, {13'sd-2162, 10'sd-475, 13'sd-2079}},
{{12'sd-1664, 12'sd-1434, 13'sd-2174}, {12'sd1305, 13'sd-2199, 12'sd-1238}, {12'sd-1274, 12'sd-1519, 11'sd586}},
{{12'sd-1065, 12'sd1962, 11'sd-815}, {13'sd-2886, 13'sd2163, 10'sd451}, {12'sd1903, 12'sd-1387, 11'sd-595}},
{{13'sd-2203, 13'sd-2081, 10'sd492}, {11'sd-689, 12'sd-1736, 13'sd2813}, {12'sd1607, 12'sd-1777, 11'sd611}},
{{13'sd-2489, 12'sd1238, 13'sd2141}, {12'sd1105, 13'sd2237, 13'sd-2708}, {13'sd-2656, 13'sd-2547, 13'sd-2422}},
{{12'sd1542, 11'sd939, 11'sd823}, {13'sd-2221, 12'sd1432, 13'sd2216}, {13'sd2413, 13'sd2581, 8'sd-112}},
{{11'sd-569, 11'sd548, 12'sd1377}, {13'sd2457, 12'sd1826, 11'sd-747}, {13'sd-2876, 12'sd1136, 12'sd1262}},
{{13'sd2189, 11'sd-858, 10'sd-307}, {11'sd-814, 13'sd2791, 12'sd1912}, {12'sd-1174, 12'sd1359, 12'sd1452}},
{{13'sd-2266, 10'sd-345, 13'sd-2551}, {13'sd-2158, 12'sd-1482, 12'sd1986}, {13'sd2963, 13'sd2283, 9'sd-186}},
{{11'sd-637, 13'sd-2196, 13'sd-2550}, {13'sd-2858, 11'sd-818, 13'sd-2690}, {13'sd-2738, 10'sd450, 12'sd1821}},
{{12'sd2041, 11'sd-772, 13'sd-2174}, {13'sd-2991, 12'sd-1876, 9'sd189}, {11'sd-988, 12'sd-1183, 13'sd-2759}},
{{11'sd-958, 13'sd2121, 10'sd-442}, {12'sd1644, 12'sd1309, 13'sd2363}, {13'sd-2340, 13'sd-2397, 13'sd-2234}},
{{11'sd-928, 13'sd-2410, 11'sd-539}, {11'sd907, 12'sd-1620, 10'sd308}, {9'sd223, 11'sd785, 12'sd1387}},
{{10'sd445, 11'sd-933, 8'sd-96}, {12'sd1179, 13'sd-2521, 10'sd-260}, {12'sd-1281, 11'sd-557, 11'sd896}},
{{13'sd-2231, 13'sd-3233, 11'sd1005}, {10'sd380, 10'sd-495, 13'sd-2170}, {11'sd548, 12'sd1159, 13'sd2228}},
{{12'sd-1111, 13'sd2832, 12'sd-1210}, {9'sd-213, 11'sd660, 12'sd1500}, {10'sd-319, 13'sd2404, 13'sd-2474}},
{{11'sd-601, 12'sd1732, 12'sd1329}, {13'sd-2628, 11'sd787, 10'sd-320}, {11'sd625, 13'sd-2274, 12'sd1776}},
{{13'sd2783, 10'sd-324, 11'sd-905}, {13'sd2364, 13'sd2212, 10'sd-256}, {12'sd-1421, 13'sd-2134, 7'sd38}},
{{12'sd1108, 12'sd1434, 11'sd512}, {13'sd-2681, 12'sd-1779, 12'sd1252}, {13'sd2193, 12'sd-1398, 12'sd-1823}},
{{3'sd-3, 13'sd2553, 12'sd-1254}, {10'sd312, 11'sd754, 12'sd1535}, {12'sd-1372, 13'sd2506, 13'sd2203}}},
{
{{13'sd2253, 13'sd2500, 10'sd-400}, {13'sd2297, 13'sd-2673, 10'sd463}, {10'sd-263, 6'sd-22, 13'sd-2283}},
{{12'sd1745, 13'sd2181, 12'sd1068}, {12'sd1624, 13'sd3005, 12'sd-1154}, {12'sd1787, 13'sd2690, 13'sd2239}},
{{13'sd3278, 9'sd-147, 12'sd-1205}, {13'sd2075, 12'sd1407, 13'sd-2456}, {13'sd-3022, 11'sd926, 8'sd-68}},
{{11'sd-569, 11'sd637, 12'sd-1346}, {12'sd-1818, 8'sd-116, 8'sd113}, {11'sd699, 11'sd-785, 13'sd2160}},
{{13'sd-3233, 11'sd-593, 12'sd-1340}, {12'sd-1942, 12'sd-1312, 12'sd-1204}, {11'sd822, 12'sd1966, 12'sd1318}},
{{11'sd956, 13'sd-2399, 10'sd-426}, {13'sd-2445, 8'sd-71, 12'sd1896}, {13'sd-3142, 13'sd-2993, 11'sd-703}},
{{12'sd-1077, 12'sd-1914, 9'sd-146}, {12'sd1720, 13'sd-2878, 13'sd-2681}, {13'sd2232, 13'sd-2182, 10'sd-350}},
{{13'sd-3776, 13'sd2236, 12'sd1722}, {12'sd1655, 13'sd2254, 13'sd3399}, {12'sd-1817, 13'sd-3082, 12'sd1117}},
{{13'sd3085, 10'sd506, 12'sd-1648}, {12'sd1993, 11'sd-908, 12'sd1285}, {11'sd-620, 12'sd1638, 12'sd1370}},
{{11'sd-782, 11'sd829, 9'sd234}, {12'sd-1982, 9'sd-183, 10'sd-511}, {11'sd-706, 13'sd2498, 12'sd-1586}},
{{6'sd-17, 13'sd-3030, 12'sd-1801}, {13'sd-2056, 12'sd1080, 12'sd1089}, {11'sd539, 13'sd3453, 14'sd5100}},
{{11'sd903, 13'sd-3058, 12'sd-1624}, {12'sd1192, 7'sd44, 11'sd-944}, {13'sd2323, 11'sd818, 7'sd-62}},
{{13'sd-3699, 13'sd-2581, 13'sd-3396}, {13'sd2118, 12'sd-1628, 9'sd163}, {12'sd1853, 13'sd-2519, 12'sd-1681}},
{{13'sd-2650, 11'sd-985, 11'sd-784}, {13'sd-2162, 10'sd309, 12'sd1173}, {12'sd1914, 12'sd1699, 13'sd3229}},
{{13'sd-2854, 11'sd1007, 11'sd-881}, {11'sd-891, 11'sd-818, 13'sd-2603}, {12'sd1422, 11'sd660, 12'sd-1204}},
{{12'sd1792, 12'sd1772, 13'sd-2129}, {12'sd1671, 13'sd2291, 11'sd838}, {13'sd2654, 11'sd-558, 12'sd1858}},
{{11'sd-816, 11'sd-593, 12'sd-1098}, {13'sd2779, 11'sd-534, 11'sd-648}, {13'sd2721, 11'sd847, 9'sd-254}},
{{12'sd1695, 12'sd-1699, 9'sd-153}, {9'sd237, 13'sd-3254, 11'sd610}, {13'sd-2093, 11'sd-565, 12'sd-1615}},
{{13'sd2585, 12'sd-1136, 12'sd1978}, {11'sd984, 12'sd1282, 7'sd-44}, {12'sd-1221, 12'sd-1279, 12'sd1416}},
{{13'sd-2458, 10'sd-378, 12'sd-1893}, {13'sd2565, 12'sd-1817, 11'sd805}, {9'sd-225, 12'sd-1478, 12'sd-1954}},
{{13'sd2873, 11'sd-928, 12'sd-1421}, {10'sd309, 13'sd-2505, 12'sd-1756}, {12'sd1809, 12'sd-1417, 12'sd1516}},
{{7'sd47, 12'sd1960, 12'sd-1274}, {12'sd1395, 13'sd-2873, 9'sd-238}, {9'sd143, 14'sd4243, 13'sd2106}},
{{13'sd3111, 11'sd-803, 11'sd966}, {12'sd1385, 12'sd1206, 11'sd649}, {11'sd838, 12'sd2001, 13'sd2273}},
{{11'sd534, 11'sd787, 12'sd-1914}, {13'sd2240, 11'sd649, 10'sd-323}, {10'sd425, 11'sd619, 12'sd1558}},
{{12'sd1356, 13'sd2423, 13'sd-2114}, {12'sd1027, 6'sd-25, 13'sd-2705}, {11'sd-1015, 9'sd-208, 13'sd-4046}},
{{13'sd-2397, 7'sd-32, 12'sd-1550}, {13'sd2112, 12'sd-1174, 13'sd2444}, {12'sd1585, 11'sd-905, 13'sd2371}},
{{12'sd1179, 3'sd3, 12'sd-1373}, {13'sd2633, 11'sd-731, 11'sd-937}, {8'sd-79, 9'sd-216, 12'sd-1058}},
{{11'sd774, 12'sd-1455, 13'sd3084}, {12'sd1423, 11'sd913, 13'sd2058}, {10'sd507, 11'sd-867, 12'sd-1230}},
{{13'sd-2343, 13'sd-3202, 12'sd-1835}, {13'sd-3052, 12'sd1937, 12'sd-1596}, {12'sd1406, 9'sd-145, 13'sd2417}},
{{14'sd-4212, 13'sd-2191, 12'sd1227}, {10'sd395, 12'sd-1815, 12'sd-1772}, {12'sd1999, 9'sd240, 13'sd3118}},
{{10'sd-498, 13'sd2573, 13'sd-2177}, {12'sd1710, 12'sd-1746, 12'sd1159}, {13'sd-2576, 12'sd-1590, 9'sd201}},
{{13'sd-2058, 12'sd1227, 12'sd1410}, {12'sd1024, 13'sd2888, 12'sd-1550}, {12'sd-1963, 12'sd-1751, 11'sd718}},
{{11'sd1004, 12'sd-1641, 13'sd-2714}, {12'sd-1710, 12'sd-1487, 13'sd-2340}, {12'sd1782, 13'sd-2783, 12'sd1643}},
{{13'sd2805, 13'sd2368, 13'sd-2151}, {13'sd-2563, 13'sd2459, 13'sd-2451}, {10'sd-459, 11'sd-531, 12'sd1767}},
{{10'sd-439, 10'sd-380, 10'sd434}, {13'sd2186, 8'sd-102, 12'sd1973}, {13'sd-2400, 11'sd-970, 11'sd871}},
{{13'sd-2226, 12'sd1355, 13'sd2317}, {11'sd-600, 9'sd247, 11'sd696}, {12'sd-1926, 10'sd-379, 12'sd-1093}},
{{12'sd-1301, 10'sd-260, 13'sd3263}, {7'sd-43, 11'sd-573, 12'sd1237}, {13'sd-2438, 13'sd-2343, 12'sd-1910}},
{{9'sd-211, 10'sd421, 13'sd-2441}, {13'sd2542, 13'sd2815, 13'sd2793}, {13'sd3773, 13'sd3523, 10'sd464}},
{{11'sd-618, 13'sd-2114, 11'sd877}, {13'sd2585, 13'sd2827, 12'sd1676}, {11'sd1000, 13'sd3440, 12'sd1934}},
{{12'sd1496, 9'sd-217, 7'sd-54}, {10'sd-340, 12'sd1478, 10'sd461}, {13'sd2692, 12'sd1786, 11'sd-917}},
{{12'sd-1570, 9'sd145, 11'sd-747}, {13'sd2451, 12'sd-1383, 12'sd-1942}, {13'sd-2271, 13'sd-2597, 12'sd-1180}},
{{12'sd1704, 12'sd-1372, 13'sd2425}, {12'sd-1332, 6'sd24, 12'sd1258}, {13'sd2461, 10'sd457, 12'sd-1038}},
{{11'sd-916, 12'sd1577, 10'sd424}, {10'sd-342, 11'sd-743, 2'sd-1}, {9'sd240, 13'sd-3037, 12'sd1796}},
{{10'sd509, 13'sd2785, 11'sd809}, {11'sd734, 12'sd1999, 13'sd2691}, {11'sd538, 7'sd-58, 11'sd-937}},
{{11'sd-575, 13'sd-2322, 12'sd-1519}, {13'sd-2725, 13'sd-2923, 13'sd2243}, {11'sd-743, 10'sd355, 11'sd-738}},
{{13'sd2538, 13'sd2965, 10'sd-424}, {12'sd-1237, 13'sd2161, 12'sd1196}, {12'sd1070, 11'sd806, 12'sd-1661}},
{{12'sd-1273, 8'sd99, 13'sd-2093}, {11'sd881, 13'sd-2687, 13'sd-3189}, {10'sd-457, 13'sd-2372, 12'sd-1992}},
{{13'sd2083, 12'sd-1625, 11'sd-710}, {13'sd-2523, 13'sd-2531, 12'sd1830}, {13'sd2494, 12'sd-1262, 13'sd2058}},
{{11'sd-958, 13'sd-2467, 13'sd-2206}, {13'sd-2925, 13'sd-2533, 12'sd-1343}, {12'sd-1843, 11'sd998, 12'sd-1999}},
{{13'sd-2873, 13'sd-2664, 5'sd-10}, {13'sd-2344, 12'sd-2026, 12'sd-1304}, {11'sd-730, 10'sd375, 12'sd1248}},
{{12'sd1329, 10'sd380, 13'sd-2580}, {13'sd-2125, 11'sd-960, 12'sd1620}, {12'sd1182, 11'sd984, 12'sd-1613}},
{{13'sd-2826, 12'sd-1064, 12'sd-1217}, {12'sd2009, 12'sd-1082, 12'sd-1482}, {12'sd1806, 11'sd-669, 13'sd2897}},
{{13'sd-2505, 13'sd-2171, 9'sd-184}, {11'sd933, 13'sd-2735, 9'sd-131}, {12'sd2036, 11'sd739, 14'sd4734}},
{{13'sd2927, 13'sd-2072, 10'sd-318}, {9'sd191, 11'sd-672, 13'sd-2520}, {11'sd-805, 13'sd-2270, 12'sd-1056}},
{{13'sd-2196, 9'sd162, 12'sd1136}, {11'sd-646, 10'sd-371, 13'sd-2610}, {12'sd1742, 10'sd261, 12'sd1428}},
{{9'sd131, 11'sd-762, 13'sd-2108}, {11'sd740, 9'sd163, 12'sd-1055}, {13'sd-2215, 13'sd-2793, 13'sd-2884}},
{{11'sd636, 12'sd-1666, 13'sd-2559}, {12'sd1631, 12'sd1799, 11'sd660}, {13'sd2491, 13'sd2103, 9'sd249}},
{{11'sd727, 11'sd-649, 13'sd2939}, {13'sd2197, 9'sd220, 12'sd-1619}, {13'sd-2059, 11'sd595, 11'sd785}},
{{12'sd1653, 11'sd-1020, 13'sd2146}, {12'sd-1572, 12'sd-1394, 12'sd1239}, {14'sd-4841, 13'sd-2826, 12'sd-1951}},
{{13'sd-2164, 11'sd941, 13'sd2395}, {11'sd866, 13'sd2170, 11'sd-741}, {10'sd-300, 10'sd-459, 11'sd-980}},
{{8'sd-80, 11'sd-782, 13'sd-2982}, {12'sd1815, 11'sd-962, 13'sd2071}, {13'sd-2761, 12'sd-1281, 12'sd-1545}},
{{13'sd-2763, 9'sd177, 8'sd-88}, {11'sd-891, 12'sd1266, 11'sd-862}, {11'sd925, 11'sd-824, 13'sd3178}},
{{12'sd1707, 8'sd98, 13'sd-2668}, {11'sd992, 11'sd969, 12'sd-1727}, {12'sd-1441, 12'sd-1036, 13'sd-2431}},
{{12'sd-1604, 12'sd-1745, 12'sd1172}, {12'sd-1965, 13'sd-2054, 12'sd-1068}, {12'sd-1382, 12'sd-2038, 13'sd2644}}},
{
{{9'sd-244, 9'sd212, 13'sd-3903}, {11'sd-946, 12'sd1695, 12'sd-1673}, {13'sd2707, 11'sd-958, 11'sd642}},
{{13'sd-2165, 9'sd-240, 11'sd-1004}, {13'sd-2279, 11'sd945, 8'sd77}, {11'sd535, 13'sd-2955, 12'sd1384}},
{{13'sd-2589, 11'sd515, 12'sd-1180}, {11'sd-872, 13'sd2343, 13'sd2065}, {9'sd-160, 12'sd1693, 12'sd1910}},
{{12'sd-1325, 12'sd2030, 11'sd-616}, {13'sd-2546, 12'sd1042, 13'sd-2201}, {11'sd-819, 12'sd1844, 11'sd-809}},
{{12'sd-1930, 11'sd-747, 10'sd448}, {11'sd804, 7'sd42, 8'sd125}, {12'sd-1375, 12'sd-2024, 9'sd-199}},
{{13'sd-2692, 11'sd-679, 12'sd-1763}, {12'sd-1331, 11'sd998, 12'sd1787}, {13'sd2712, 13'sd2767, 10'sd422}},
{{12'sd1201, 12'sd-1605, 12'sd1640}, {11'sd927, 12'sd-1626, 8'sd71}, {13'sd2122, 11'sd738, 14'sd-4198}},
{{12'sd-1929, 11'sd981, 11'sd-556}, {6'sd20, 12'sd1980, 14'sd-4169}, {11'sd591, 12'sd-1148, 13'sd-3517}},
{{13'sd-2638, 11'sd-531, 13'sd2153}, {12'sd1279, 12'sd1033, 11'sd-720}, {10'sd-383, 12'sd1817, 9'sd-190}},
{{12'sd1250, 12'sd1221, 12'sd1840}, {12'sd1604, 12'sd-1302, 11'sd-860}, {12'sd-1205, 12'sd1333, 10'sd-262}},
{{13'sd2065, 12'sd1687, 13'sd-2091}, {13'sd-2107, 10'sd-372, 13'sd-2891}, {9'sd-173, 13'sd-2080, 13'sd-2877}},
{{13'sd-3067, 12'sd1903, 11'sd863}, {11'sd572, 12'sd1280, 13'sd-2427}, {13'sd2539, 13'sd2972, 13'sd-2409}},
{{11'sd946, 12'sd1803, 13'sd3181}, {12'sd-2034, 7'sd-58, 12'sd1652}, {10'sd-467, 12'sd-1063, 11'sd-757}},
{{11'sd-893, 12'sd1496, 12'sd-1262}, {12'sd1638, 13'sd-2242, 12'sd-1214}, {13'sd2300, 11'sd-822, 12'sd-1619}},
{{10'sd-437, 13'sd2980, 13'sd2357}, {13'sd2300, 11'sd838, 12'sd1515}, {12'sd1355, 12'sd-1435, 11'sd639}},
{{10'sd301, 12'sd-1380, 10'sd-503}, {13'sd-2112, 12'sd1982, 12'sd-1566}, {12'sd-1317, 13'sd-2758, 13'sd-3094}},
{{9'sd-212, 12'sd-1957, 7'sd-56}, {13'sd-2306, 12'sd1172, 11'sd975}, {13'sd-2063, 8'sd68, 11'sd796}},
{{10'sd-386, 13'sd2358, 14'sd4656}, {8'sd88, 14'sd-4141, 11'sd-760}, {13'sd4018, 12'sd-1860, 13'sd2197}},
{{12'sd1403, 9'sd208, 9'sd-229}, {12'sd1874, 13'sd2103, 7'sd-37}, {12'sd-2028, 11'sd713, 13'sd-2092}},
{{11'sd885, 9'sd218, 11'sd541}, {8'sd113, 11'sd-871, 13'sd3201}, {12'sd1581, 12'sd-1436, 11'sd989}},
{{11'sd890, 11'sd-634, 12'sd-1122}, {13'sd-2210, 12'sd-1178, 13'sd3688}, {13'sd2373, 12'sd-1553, 13'sd2304}},
{{12'sd-1396, 13'sd3510, 8'sd-87}, {10'sd-498, 12'sd-1173, 13'sd-2400}, {12'sd-1666, 13'sd-3015, 11'sd-720}},
{{11'sd-960, 11'sd-592, 13'sd2495}, {12'sd-1250, 13'sd2272, 9'sd-193}, {12'sd-1344, 13'sd-2843, 10'sd261}},
{{11'sd-575, 12'sd-1516, 11'sd655}, {12'sd-1831, 11'sd-617, 13'sd2623}, {12'sd1863, 12'sd-1951, 9'sd247}},
{{11'sd739, 13'sd-3302, 13'sd-2881}, {9'sd166, 13'sd2236, 13'sd2673}, {11'sd781, 13'sd2864, 13'sd3847}},
{{12'sd-1505, 13'sd-2414, 12'sd-1775}, {12'sd1254, 12'sd-1920, 12'sd-1665}, {9'sd-185, 12'sd1198, 10'sd-449}},
{{13'sd2128, 11'sd533, 13'sd-2802}, {12'sd-1400, 13'sd2110, 11'sd554}, {13'sd2265, 11'sd-803, 9'sd-172}},
{{10'sd-295, 12'sd1818, 12'sd1081}, {11'sd1000, 13'sd-2867, 11'sd772}, {11'sd-746, 13'sd2765, 12'sd1547}},
{{12'sd-1544, 13'sd2915, 13'sd2381}, {12'sd1474, 12'sd1959, 12'sd-1780}, {13'sd-2554, 13'sd-3050, 12'sd1149}},
{{13'sd3387, 12'sd-1291, 13'sd-2795}, {13'sd2051, 12'sd1042, 11'sd-524}, {11'sd-621, 13'sd-2312, 11'sd-732}},
{{12'sd1954, 12'sd1876, 11'sd-555}, {11'sd-978, 13'sd2819, 13'sd2785}, {13'sd-2844, 6'sd-26, 13'sd-2262}},
{{12'sd-1935, 10'sd-503, 13'sd-2109}, {13'sd-2422, 12'sd-1659, 12'sd-1064}, {12'sd-1444, 12'sd1320, 13'sd-2489}},
{{12'sd1293, 12'sd-1233, 13'sd2519}, {11'sd-965, 12'sd1141, 13'sd-2086}, {12'sd-1947, 13'sd-2753, 11'sd548}},
{{11'sd-997, 10'sd-318, 13'sd2314}, {12'sd1114, 12'sd1794, 11'sd584}, {12'sd-1377, 12'sd-1981, 13'sd3573}},
{{9'sd-199, 12'sd-1473, 14'sd-4289}, {11'sd-929, 11'sd-704, 13'sd-3699}, {13'sd3382, 11'sd565, 12'sd1300}},
{{12'sd-1713, 12'sd1996, 11'sd692}, {13'sd2100, 12'sd-1436, 10'sd411}, {12'sd-1079, 13'sd2152, 11'sd-883}},
{{11'sd559, 11'sd-973, 13'sd2834}, {11'sd-903, 13'sd2551, 13'sd2569}, {11'sd-543, 13'sd-2892, 13'sd-2119}},
{{10'sd294, 10'sd378, 12'sd-1137}, {9'sd-148, 10'sd-319, 12'sd-1428}, {12'sd1424, 13'sd-3607, 14'sd-4508}},
{{11'sd-986, 10'sd374, 10'sd299}, {12'sd-1859, 11'sd-850, 10'sd-403}, {13'sd-3546, 13'sd-3268, 13'sd-3203}},
{{13'sd2268, 12'sd1598, 12'sd1646}, {13'sd-3050, 8'sd-116, 13'sd-3079}, {10'sd-392, 11'sd993, 11'sd1003}},
{{12'sd-1331, 13'sd-2775, 12'sd-1290}, {13'sd-2327, 12'sd1181, 7'sd50}, {12'sd-1396, 12'sd-1256, 13'sd2707}},
{{9'sd-163, 12'sd1671, 9'sd-237}, {10'sd-383, 10'sd-338, 12'sd-1300}, {12'sd-1172, 11'sd-666, 13'sd2679}},
{{10'sd279, 13'sd2140, 12'sd1809}, {12'sd-1540, 11'sd-778, 7'sd-39}, {13'sd2602, 13'sd3148, 13'sd-2343}},
{{13'sd-2191, 10'sd-389, 12'sd-1465}, {10'sd-341, 13'sd2625, 12'sd-1716}, {9'sd-247, 12'sd1205, 13'sd3254}},
{{13'sd2488, 11'sd-559, 12'sd1167}, {11'sd-525, 11'sd-723, 12'sd-1110}, {12'sd1823, 8'sd-67, 11'sd554}},
{{12'sd-1077, 12'sd1166, 13'sd2339}, {11'sd894, 12'sd1716, 11'sd-605}, {11'sd-851, 12'sd-1307, 10'sd-326}},
{{8'sd78, 12'sd-1993, 12'sd1221}, {12'sd-1708, 13'sd-3274, 13'sd-2317}, {12'sd1436, 13'sd-3369, 12'sd1985}},
{{13'sd-2073, 13'sd2327, 11'sd-1003}, {11'sd-728, 12'sd-1896, 13'sd2124}, {13'sd-2427, 12'sd1700, 11'sd926}},
{{12'sd1710, 11'sd-986, 9'sd-245}, {12'sd-1841, 12'sd-1707, 11'sd645}, {7'sd58, 13'sd3215, 13'sd2402}},
{{12'sd-1676, 12'sd1740, 11'sd726}, {9'sd128, 11'sd615, 13'sd2338}, {7'sd47, 13'sd-2627, 10'sd421}},
{{12'sd1257, 10'sd434, 13'sd2290}, {11'sd843, 12'sd-1399, 13'sd-2698}, {9'sd178, 13'sd-2257, 12'sd-1682}},
{{12'sd-1948, 13'sd2336, 12'sd1685}, {12'sd1966, 13'sd2057, 13'sd-2749}, {13'sd2232, 13'sd-2196, 10'sd-382}},
{{11'sd582, 13'sd4090, 13'sd3467}, {9'sd241, 12'sd-1373, 11'sd-609}, {11'sd900, 12'sd-1867, 12'sd-1777}},
{{11'sd-646, 12'sd-1105, 10'sd272}, {12'sd1075, 9'sd-245, 13'sd-2438}, {13'sd-2411, 11'sd-521, 12'sd1590}},
{{12'sd-1288, 8'sd108, 13'sd-2049}, {13'sd-2185, 8'sd-91, 12'sd1525}, {9'sd154, 10'sd428, 13'sd-2101}},
{{12'sd-1429, 11'sd514, 12'sd-1856}, {12'sd1086, 6'sd-24, 12'sd-1762}, {12'sd-1072, 12'sd1804, 11'sd794}},
{{13'sd2274, 10'sd385, 13'sd2702}, {12'sd1804, 11'sd837, 12'sd-1336}, {13'sd-2530, 12'sd-1314, 12'sd1865}},
{{13'sd-2289, 11'sd949, 12'sd-1873}, {12'sd1523, 11'sd-841, 13'sd-3803}, {11'sd-584, 13'sd2749, 11'sd810}},
{{13'sd-2115, 13'sd-2976, 12'sd-1625}, {13'sd2618, 12'sd1096, 13'sd-2904}, {14'sd6409, 13'sd2684, 12'sd1827}},
{{10'sd511, 13'sd-2619, 12'sd-1058}, {11'sd517, 10'sd-460, 9'sd228}, {12'sd-2008, 13'sd2599, 12'sd-1105}},
{{11'sd759, 13'sd-2718, 10'sd-374}, {12'sd-1595, 11'sd-834, 12'sd-1448}, {12'sd1663, 13'sd3127, 13'sd2133}},
{{12'sd1618, 12'sd2044, 13'sd-2676}, {12'sd-1071, 13'sd-2346, 11'sd748}, {10'sd-339, 7'sd-54, 12'sd-1046}},
{{10'sd505, 7'sd54, 13'sd3438}, {5'sd-12, 12'sd-1035, 14'sd4644}, {12'sd1336, 12'sd1541, 11'sd-561}},
{{13'sd-2670, 12'sd-1081, 11'sd-895}, {13'sd2172, 13'sd2114, 11'sd730}, {13'sd-2658, 12'sd-1263, 13'sd-2076}}},
{
{{13'sd-2364, 11'sd-666, 8'sd68}, {10'sd448, 13'sd-2120, 12'sd-1409}, {12'sd1586, 10'sd340, 10'sd-336}},
{{11'sd642, 10'sd-483, 12'sd-1134}, {12'sd1369, 9'sd-230, 8'sd92}, {12'sd-1717, 13'sd2616, 12'sd1984}},
{{11'sd615, 13'sd2203, 13'sd-2987}, {8'sd92, 11'sd-942, 13'sd-2765}, {12'sd-1615, 10'sd-293, 10'sd279}},
{{12'sd-2037, 11'sd-580, 12'sd-1884}, {10'sd415, 13'sd-3086, 13'sd-2633}, {10'sd367, 12'sd-1763, 11'sd824}},
{{12'sd1466, 12'sd-1480, 11'sd1019}, {12'sd-1052, 8'sd100, 7'sd-55}, {11'sd-570, 10'sd-282, 12'sd1852}},
{{13'sd2768, 13'sd2572, 9'sd202}, {13'sd-2942, 12'sd1604, 11'sd-530}, {12'sd-1795, 13'sd2444, 12'sd-1646}},
{{13'sd2526, 10'sd274, 13'sd2389}, {10'sd422, 13'sd-2451, 12'sd-1232}, {13'sd2144, 13'sd-2710, 11'sd681}},
{{12'sd1216, 12'sd-1513, 11'sd-789}, {13'sd-2250, 12'sd-1557, 11'sd676}, {11'sd816, 11'sd973, 12'sd-1280}},
{{11'sd-877, 12'sd-1603, 13'sd-2066}, {12'sd1604, 13'sd2390, 11'sd582}, {11'sd-528, 11'sd879, 11'sd-528}},
{{11'sd-519, 8'sd109, 9'sd-137}, {12'sd-1471, 12'sd1289, 13'sd3115}, {13'sd2659, 11'sd-996, 12'sd1762}},
{{12'sd-1643, 10'sd-357, 12'sd1956}, {12'sd-1287, 13'sd-2269, 12'sd1834}, {14'sd-5037, 14'sd-5363, 12'sd1971}},
{{13'sd2305, 11'sd-642, 12'sd-1855}, {11'sd-926, 12'sd1854, 11'sd830}, {12'sd1649, 8'sd70, 11'sd-967}},
{{13'sd2161, 13'sd-2392, 13'sd-3108}, {13'sd3031, 12'sd-1300, 11'sd-716}, {10'sd-405, 12'sd1406, 11'sd778}},
{{10'sd-273, 13'sd2071, 12'sd1099}, {12'sd-1894, 5'sd8, 11'sd-1003}, {12'sd1889, 11'sd801, 12'sd-1969}},
{{12'sd-2022, 9'sd135, 11'sd-810}, {12'sd-1312, 6'sd26, 13'sd2416}, {12'sd1459, 12'sd1894, 12'sd1737}},
{{12'sd-1867, 12'sd1396, 13'sd2201}, {11'sd-570, 13'sd-2398, 10'sd-349}, {13'sd2861, 11'sd-938, 12'sd1985}},
{{13'sd2388, 13'sd-2472, 13'sd2238}, {11'sd591, 12'sd-1730, 8'sd-122}, {13'sd3111, 11'sd653, 12'sd-1174}},
{{12'sd-1802, 9'sd156, 12'sd1104}, {12'sd1559, 11'sd-906, 8'sd123}, {13'sd4083, 11'sd765, 13'sd3089}},
{{5'sd-9, 11'sd946, 11'sd932}, {12'sd-1154, 11'sd-891, 13'sd-2244}, {11'sd-675, 11'sd538, 12'sd-1416}},
{{13'sd2212, 13'sd-2777, 9'sd227}, {10'sd317, 12'sd1172, 13'sd-2137}, {11'sd-750, 12'sd-2023, 13'sd2080}},
{{13'sd2606, 12'sd-1749, 13'sd-2083}, {11'sd572, 12'sd1087, 11'sd-920}, {13'sd-2632, 13'sd2173, 13'sd2219}},
{{12'sd1591, 11'sd-932, 11'sd702}, {11'sd-695, 13'sd-2521, 9'sd154}, {8'sd110, 12'sd-1724, 12'sd1541}},
{{12'sd-1586, 12'sd1514, 7'sd62}, {12'sd-1883, 11'sd1000, 9'sd139}, {12'sd-1979, 4'sd4, 12'sd-1458}},
{{12'sd-1967, 11'sd-549, 12'sd1846}, {13'sd-2548, 12'sd1569, 12'sd-1846}, {12'sd-1276, 11'sd624, 11'sd-823}},
{{13'sd2918, 12'sd1400, 12'sd1637}, {12'sd1362, 12'sd-1028, 11'sd-836}, {12'sd1709, 14'sd4773, 10'sd-311}},
{{12'sd-1659, 9'sd249, 12'sd-1592}, {10'sd341, 13'sd2724, 11'sd659}, {12'sd-1155, 13'sd-2211, 12'sd1729}},
{{12'sd1758, 11'sd-957, 13'sd-2093}, {11'sd-798, 12'sd-1986, 13'sd-2474}, {12'sd-1145, 12'sd1666, 9'sd177}},
{{11'sd1007, 13'sd2456, 10'sd-407}, {12'sd1679, 13'sd2881, 11'sd694}, {12'sd1113, 10'sd504, 12'sd1749}},
{{12'sd-1672, 11'sd-718, 12'sd1456}, {12'sd1290, 10'sd318, 9'sd-193}, {11'sd719, 10'sd325, 13'sd2078}},
{{11'sd-619, 13'sd-2543, 12'sd-1478}, {10'sd-287, 12'sd1699, 6'sd30}, {11'sd519, 12'sd1832, 12'sd1524}},
{{13'sd-2937, 12'sd1166, 13'sd2289}, {11'sd-900, 8'sd94, 13'sd-2443}, {11'sd638, 11'sd-1008, 11'sd984}},
{{10'sd-510, 13'sd2157, 12'sd2047}, {12'sd1973, 11'sd866, 11'sd-974}, {8'sd113, 13'sd2621, 12'sd-1986}},
{{13'sd2234, 11'sd665, 9'sd146}, {8'sd-117, 12'sd-1812, 13'sd2538}, {12'sd-1661, 12'sd1817, 12'sd1492}},
{{9'sd164, 13'sd2845, 12'sd-1999}, {12'sd1775, 10'sd-465, 10'sd463}, {10'sd325, 13'sd-2638, 13'sd-2262}},
{{13'sd2221, 13'sd-2481, 8'sd123}, {11'sd977, 8'sd-91, 11'sd957}, {10'sd337, 10'sd312, 12'sd1140}},
{{13'sd2375, 12'sd-1692, 12'sd-1688}, {13'sd-2662, 7'sd-59, 12'sd1907}, {12'sd-1560, 12'sd-1629, 10'sd321}},
{{11'sd-575, 11'sd695, 11'sd643}, {11'sd536, 12'sd-1380, 13'sd2282}, {13'sd-3344, 11'sd714, 12'sd-1167}},
{{12'sd-1303, 11'sd-805, 13'sd-2662}, {13'sd-2666, 12'sd1376, 12'sd1753}, {12'sd1980, 13'sd2904, 12'sd-1570}},
{{13'sd2330, 11'sd-815, 12'sd-1497}, {11'sd-818, 13'sd-3114, 11'sd992}, {13'sd2625, 12'sd-1602, 13'sd-2776}},
{{10'sd274, 12'sd-1977, 12'sd1885}, {11'sd948, 13'sd-2807, 12'sd1328}, {13'sd2340, 11'sd551, 11'sd-734}},
{{8'sd-107, 13'sd2143, 13'sd-2348}, {11'sd527, 12'sd-1727, 12'sd-1437}, {10'sd-343, 13'sd-2176, 13'sd-2128}},
{{12'sd1763, 11'sd608, 12'sd1703}, {12'sd-1559, 9'sd-156, 12'sd-1500}, {11'sd597, 13'sd-2094, 13'sd2302}},
{{11'sd792, 12'sd-1277, 12'sd-1397}, {11'sd-927, 6'sd29, 12'sd2045}, {12'sd1038, 11'sd985, 11'sd952}},
{{11'sd740, 13'sd2619, 12'sd1662}, {11'sd-963, 7'sd36, 13'sd-3203}, {11'sd997, 12'sd1236, 12'sd-2039}},
{{13'sd-2195, 12'sd1139, 12'sd-1870}, {12'sd1292, 12'sd1745, 12'sd-1189}, {13'sd-2920, 12'sd-1781, 13'sd2475}},
{{12'sd-1034, 12'sd-1553, 10'sd-403}, {10'sd-275, 12'sd1656, 11'sd-962}, {9'sd-196, 13'sd2108, 12'sd1880}},
{{12'sd1537, 12'sd1306, 12'sd-1749}, {12'sd1372, 12'sd-1360, 11'sd-996}, {11'sd-576, 12'sd1796, 12'sd-1865}},
{{12'sd1066, 13'sd2059, 12'sd1801}, {11'sd859, 8'sd-104, 12'sd-1790}, {12'sd1572, 10'sd-430, 12'sd-1733}},
{{13'sd2451, 10'sd-328, 11'sd-585}, {13'sd-2214, 13'sd-2170, 12'sd-1180}, {12'sd-1389, 12'sd1361, 13'sd2408}},
{{12'sd-1689, 10'sd-269, 13'sd-2589}, {12'sd1499, 11'sd-518, 13'sd2140}, {12'sd-1747, 12'sd1965, 13'sd2192}},
{{9'sd-217, 11'sd-1016, 12'sd-1046}, {13'sd-2121, 13'sd2319, 12'sd1679}, {9'sd-198, 12'sd-1533, 12'sd-1849}},
{{13'sd-2399, 12'sd1741, 12'sd1159}, {12'sd-1664, 13'sd2547, 12'sd-1959}, {13'sd2421, 9'sd217, 11'sd741}},
{{13'sd2433, 11'sd724, 10'sd-499}, {9'sd-243, 12'sd-1030, 10'sd390}, {12'sd-1236, 13'sd2218, 10'sd260}},
{{13'sd-2637, 10'sd487, 13'sd-2172}, {12'sd1137, 12'sd1229, 12'sd1793}, {13'sd-2292, 12'sd-1987, 7'sd-50}},
{{11'sd-767, 11'sd647, 12'sd1371}, {13'sd-2224, 12'sd-1122, 13'sd-2217}, {13'sd-2588, 13'sd2412, 11'sd589}},
{{13'sd-2728, 13'sd2298, 9'sd242}, {13'sd-2280, 13'sd3010, 12'sd1148}, {12'sd-1748, 12'sd1895, 13'sd2229}},
{{12'sd1181, 11'sd868, 7'sd-46}, {10'sd328, 13'sd2640, 10'sd384}, {12'sd-1036, 12'sd1778, 11'sd-979}},
{{11'sd-803, 11'sd681, 13'sd2779}, {13'sd3096, 13'sd2637, 10'sd-404}, {13'sd3892, 9'sd-165, 12'sd-1440}},
{{10'sd334, 13'sd2488, 12'sd1584}, {12'sd-1326, 13'sd2281, 13'sd2127}, {13'sd2569, 12'sd-1252, 13'sd-3570}},
{{11'sd920, 12'sd-1536, 13'sd-2223}, {8'sd97, 12'sd1397, 13'sd-2161}, {11'sd-908, 9'sd238, 12'sd1996}},
{{11'sd-1006, 11'sd-905, 11'sd-551}, {11'sd-722, 13'sd2714, 9'sd-206}, {11'sd621, 10'sd-382, 12'sd-1698}},
{{13'sd-2509, 12'sd1209, 13'sd-2167}, {13'sd2135, 11'sd-941, 12'sd1129}, {13'sd2066, 13'sd2703, 13'sd2840}},
{{11'sd-623, 10'sd424, 10'sd-495}, {13'sd-2053, 13'sd2101, 13'sd-2629}, {12'sd-1708, 11'sd-514, 13'sd-2238}},
{{12'sd-1252, 12'sd-1911, 13'sd2914}, {13'sd2282, 11'sd983, 11'sd-516}, {12'sd1175, 12'sd-1334, 9'sd-158}}},
{
{{13'sd3282, 12'sd1481, 13'sd2123}, {11'sd-951, 10'sd454, 12'sd1675}, {13'sd-3119, 12'sd1903, 12'sd-1449}},
{{13'sd-2223, 11'sd-769, 12'sd1534}, {12'sd1111, 12'sd1958, 11'sd735}, {12'sd-1869, 11'sd-839, 11'sd674}},
{{12'sd1968, 12'sd-1620, 12'sd-2017}, {12'sd-1873, 13'sd2310, 13'sd-3162}, {12'sd-2025, 12'sd1746, 12'sd1323}},
{{11'sd588, 13'sd-2711, 12'sd1148}, {11'sd-604, 13'sd-2418, 13'sd-2961}, {10'sd-301, 12'sd-1542, 11'sd586}},
{{12'sd1522, 12'sd1735, 13'sd3042}, {13'sd-2332, 8'sd-68, 13'sd-2051}, {12'sd-1179, 12'sd1155, 12'sd-1665}},
{{13'sd-2732, 10'sd455, 11'sd876}, {13'sd2562, 10'sd330, 10'sd381}, {13'sd-2484, 12'sd1714, 11'sd-540}},
{{11'sd968, 5'sd9, 13'sd-2544}, {9'sd133, 11'sd560, 11'sd828}, {10'sd-280, 12'sd1754, 9'sd235}},
{{12'sd-1464, 12'sd-1672, 12'sd-1415}, {12'sd1285, 10'sd-353, 13'sd-3403}, {13'sd2943, 11'sd-515, 7'sd54}},
{{10'sd-490, 12'sd1373, 13'sd-2822}, {13'sd-2270, 11'sd946, 7'sd61}, {13'sd2162, 12'sd1286, 12'sd1154}},
{{11'sd910, 11'sd573, 11'sd-649}, {12'sd-1886, 11'sd968, 13'sd-2266}, {12'sd-1401, 13'sd-2331, 11'sd579}},
{{13'sd-3116, 13'sd-3240, 11'sd-594}, {13'sd-2518, 12'sd-1702, 12'sd1273}, {11'sd816, 13'sd2592, 7'sd-38}},
{{12'sd-1112, 13'sd2260, 11'sd653}, {12'sd1659, 11'sd875, 12'sd2025}, {12'sd-1981, 11'sd-878, 11'sd-698}},
{{12'sd-1792, 9'sd212, 9'sd189}, {11'sd809, 12'sd1111, 13'sd-3239}, {13'sd2280, 12'sd-1314, 12'sd1567}},
{{11'sd706, 12'sd-1148, 13'sd2552}, {12'sd-1064, 13'sd-2778, 11'sd683}, {11'sd-1016, 9'sd-173, 11'sd-947}},
{{12'sd1493, 12'sd1066, 12'sd1150}, {12'sd1773, 10'sd278, 12'sd-1236}, {11'sd747, 12'sd-1266, 12'sd1712}},
{{12'sd2025, 12'sd1687, 10'sd460}, {9'sd243, 12'sd1233, 8'sd114}, {11'sd-750, 13'sd2208, 13'sd-2260}},
{{12'sd1880, 11'sd-819, 8'sd-98}, {13'sd3111, 13'sd2133, 12'sd-1917}, {10'sd-297, 12'sd-1766, 13'sd2134}},
{{14'sd5065, 13'sd3925, 10'sd259}, {9'sd157, 10'sd438, 13'sd-2919}, {12'sd-1100, 9'sd-248, 12'sd-1566}},
{{13'sd2378, 13'sd2426, 12'sd1796}, {13'sd2062, 11'sd-615, 12'sd-1198}, {13'sd2942, 11'sd-514, 8'sd-68}},
{{12'sd1141, 13'sd-2695, 9'sd168}, {9'sd-136, 10'sd-423, 8'sd-86}, {12'sd-1434, 12'sd1334, 13'sd2421}},
{{13'sd-2098, 3'sd-2, 10'sd-372}, {12'sd-1622, 12'sd1368, 10'sd383}, {12'sd1646, 10'sd429, 10'sd-498}},
{{9'sd196, 13'sd2167, 13'sd2127}, {13'sd-3113, 10'sd-310, 9'sd-247}, {13'sd-2426, 11'sd-839, 12'sd-1055}},
{{8'sd-111, 10'sd-428, 13'sd-2179}, {11'sd1018, 12'sd-1441, 13'sd2672}, {13'sd-2186, 12'sd1439, 9'sd163}},
{{12'sd-1611, 12'sd-1933, 12'sd-1074}, {13'sd-2635, 11'sd536, 13'sd2747}, {12'sd1487, 13'sd2247, 13'sd2549}},
{{11'sd542, 12'sd1788, 13'sd-3095}, {9'sd129, 13'sd2378, 11'sd-657}, {12'sd-1700, 12'sd1734, 12'sd1416}},
{{12'sd-1712, 11'sd906, 12'sd-1871}, {12'sd-1648, 12'sd-1439, 12'sd1113}, {13'sd2463, 10'sd-496, 12'sd1899}},
{{12'sd1128, 12'sd-1188, 12'sd1172}, {13'sd2234, 8'sd-113, 7'sd42}, {12'sd-1456, 10'sd276, 10'sd319}},
{{12'sd1525, 13'sd2336, 12'sd2013}, {13'sd2867, 9'sd-219, 12'sd-1289}, {13'sd2821, 12'sd-2024, 12'sd-1247}},
{{13'sd-2401, 12'sd1451, 12'sd1216}, {11'sd537, 12'sd-1848, 11'sd-798}, {7'sd-33, 12'sd1692, 12'sd1374}},
{{13'sd2298, 8'sd-88, 12'sd1519}, {9'sd187, 12'sd-2015, 12'sd1714}, {12'sd-1638, 12'sd-1599, 13'sd2217}},
{{13'sd-2887, 8'sd-126, 13'sd-2532}, {12'sd-1968, 11'sd861, 11'sd-586}, {13'sd-2173, 13'sd2155, 11'sd906}},
{{13'sd2314, 9'sd173, 13'sd2416}, {12'sd1440, 5'sd12, 12'sd1947}, {8'sd74, 10'sd489, 12'sd-1394}},
{{12'sd-2011, 13'sd2255, 5'sd10}, {10'sd429, 13'sd2845, 12'sd-1592}, {10'sd314, 13'sd-2269, 12'sd-1750}},
{{12'sd1393, 11'sd1022, 11'sd-908}, {10'sd419, 12'sd-1478, 10'sd-279}, {13'sd2091, 13'sd-2303, 11'sd845}},
{{11'sd593, 12'sd-1365, 13'sd-2154}, {12'sd-1343, 11'sd-988, 12'sd1990}, {12'sd-1787, 13'sd2739, 12'sd-1476}},
{{11'sd-521, 11'sd605, 11'sd-847}, {11'sd824, 13'sd-2526, 13'sd-2924}, {12'sd-1329, 12'sd-1746, 13'sd-2217}},
{{12'sd-1269, 10'sd446, 12'sd-2021}, {12'sd-1905, 11'sd-690, 12'sd-1701}, {11'sd701, 12'sd1404, 2'sd-1}},
{{12'sd1111, 10'sd432, 12'sd1025}, {8'sd-76, 11'sd749, 12'sd1278}, {12'sd-1756, 9'sd207, 13'sd-2926}},
{{12'sd1218, 11'sd-693, 13'sd-2508}, {12'sd1136, 12'sd-1087, 11'sd739}, {11'sd712, 13'sd2453, 10'sd497}},
{{11'sd-593, 13'sd2118, 10'sd385}, {11'sd-629, 13'sd-2176, 12'sd1240}, {13'sd2388, 11'sd-608, 10'sd-482}},
{{11'sd-791, 8'sd-126, 11'sd-697}, {13'sd2397, 13'sd-2448, 12'sd1956}, {12'sd1511, 11'sd650, 11'sd-606}},
{{11'sd-518, 11'sd-920, 12'sd1271}, {11'sd649, 13'sd-2673, 10'sd427}, {9'sd165, 11'sd953, 11'sd516}},
{{13'sd2266, 13'sd-2553, 13'sd2409}, {12'sd-1042, 13'sd-2454, 13'sd2130}, {10'sd328, 9'sd137, 12'sd1974}},
{{12'sd1477, 11'sd522, 11'sd-769}, {13'sd-2185, 8'sd64, 12'sd-1027}, {10'sd-475, 12'sd-1851, 13'sd2434}},
{{12'sd1344, 12'sd1323, 13'sd-2355}, {13'sd-2494, 12'sd1028, 7'sd-42}, {12'sd-1929, 12'sd-1195, 11'sd981}},
{{10'sd-421, 11'sd783, 12'sd1448}, {10'sd348, 13'sd-2502, 11'sd591}, {10'sd424, 10'sd287, 12'sd1891}},
{{12'sd-1515, 13'sd2772, 13'sd2466}, {11'sd-893, 12'sd-1471, 13'sd2444}, {12'sd-1614, 4'sd-6, 11'sd-830}},
{{12'sd-1137, 12'sd-1311, 12'sd-1329}, {12'sd1065, 13'sd2614, 12'sd1875}, {13'sd2150, 10'sd467, 12'sd-1504}},
{{13'sd2755, 13'sd-2361, 13'sd2495}, {7'sd-63, 13'sd-2827, 11'sd-741}, {10'sd-456, 12'sd-1900, 10'sd-394}},
{{11'sd996, 7'sd-52, 13'sd2546}, {12'sd-1078, 11'sd-865, 12'sd-1534}, {9'sd167, 10'sd-384, 10'sd410}},
{{9'sd-241, 12'sd1820, 9'sd-134}, {13'sd-2336, 11'sd-619, 12'sd1364}, {13'sd-2346, 12'sd1923, 12'sd1963}},
{{13'sd2720, 13'sd2209, 13'sd2654}, {11'sd-739, 11'sd-930, 12'sd-1557}, {9'sd-221, 12'sd1291, 10'sd-446}},
{{11'sd-881, 12'sd-1046, 10'sd-433}, {12'sd-1788, 11'sd820, 4'sd-6}, {12'sd1641, 12'sd1111, 12'sd-1298}},
{{12'sd-1783, 11'sd1007, 13'sd2288}, {13'sd2707, 11'sd-604, 13'sd-2158}, {11'sd-893, 13'sd-2156, 12'sd-1949}},
{{12'sd1043, 12'sd-1528, 13'sd2935}, {10'sd398, 11'sd-635, 11'sd-618}, {12'sd1171, 11'sd-787, 13'sd2254}},
{{10'sd293, 13'sd-2424, 13'sd2666}, {9'sd229, 11'sd-842, 11'sd528}, {12'sd-1322, 7'sd46, 9'sd-235}},
{{13'sd-2206, 11'sd643, 12'sd1499}, {12'sd1319, 11'sd621, 10'sd-402}, {11'sd1023, 13'sd2499, 13'sd-2644}},
{{12'sd2045, 10'sd-496, 13'sd2934}, {10'sd-448, 11'sd818, 8'sd88}, {13'sd-2626, 13'sd-2286, 13'sd-2529}},
{{10'sd-344, 10'sd354, 13'sd-2241}, {13'sd-2181, 12'sd1165, 13'sd-2231}, {13'sd-2297, 10'sd-427, 13'sd-2134}},
{{11'sd-969, 12'sd-1896, 11'sd-700}, {11'sd-712, 12'sd2028, 12'sd1523}, {11'sd-686, 11'sd-978, 8'sd85}},
{{13'sd2306, 13'sd-2622, 11'sd-652}, {10'sd471, 11'sd-985, 12'sd1840}, {12'sd1198, 9'sd-219, 10'sd-467}},
{{11'sd-603, 13'sd-2101, 12'sd-1908}, {12'sd-1662, 11'sd796, 13'sd-2051}, {13'sd2883, 11'sd694, 10'sd412}},
{{11'sd807, 13'sd-2454, 12'sd-1440}, {12'sd-1648, 13'sd2564, 11'sd-651}, {10'sd-402, 8'sd96, 12'sd1027}},
{{11'sd-726, 13'sd-2350, 13'sd2972}, {12'sd-1273, 13'sd-2091, 12'sd1448}, {12'sd1679, 12'sd-1837, 12'sd-1818}}},
{
{{12'sd1133, 12'sd1131, 12'sd1384}, {10'sd-259, 3'sd3, 9'sd-146}, {13'sd-2710, 11'sd707, 10'sd-404}},
{{9'sd254, 11'sd706, 12'sd-1762}, {9'sd-197, 11'sd710, 10'sd-374}, {11'sd658, 12'sd1027, 11'sd-783}},
{{13'sd-2825, 13'sd-2100, 13'sd-2731}, {11'sd814, 12'sd1731, 12'sd-1885}, {13'sd2700, 12'sd-1963, 12'sd1264}},
{{13'sd3152, 12'sd-1646, 13'sd2894}, {12'sd-1225, 8'sd-85, 11'sd-784}, {12'sd-1486, 12'sd1996, 10'sd282}},
{{12'sd1443, 12'sd1577, 13'sd2453}, {12'sd1555, 13'sd2114, 12'sd1189}, {12'sd1811, 11'sd-916, 10'sd-265}},
{{12'sd1559, 10'sd292, 13'sd2574}, {12'sd-1065, 11'sd753, 13'sd-2313}, {13'sd-2102, 9'sd-226, 13'sd-2430}},
{{11'sd-728, 12'sd-1092, 10'sd284}, {11'sd609, 11'sd-918, 13'sd2612}, {12'sd-1890, 12'sd-1227, 9'sd-134}},
{{12'sd1872, 11'sd712, 13'sd2052}, {13'sd2539, 11'sd615, 12'sd1965}, {12'sd1997, 13'sd-2675, 13'sd2601}},
{{10'sd-396, 9'sd166, 12'sd-2025}, {9'sd-150, 12'sd-1599, 7'sd40}, {13'sd2915, 11'sd837, 11'sd950}},
{{11'sd940, 12'sd1300, 13'sd-2082}, {12'sd1529, 10'sd-440, 13'sd-2655}, {12'sd-1487, 13'sd-2669, 10'sd439}},
{{12'sd1376, 12'sd1150, 10'sd380}, {11'sd-847, 11'sd-622, 10'sd481}, {10'sd469, 9'sd206, 8'sd-115}},
{{10'sd444, 13'sd-2241, 12'sd1244}, {10'sd-498, 11'sd918, 9'sd-247}, {12'sd1163, 12'sd-1566, 9'sd-254}},
{{12'sd1034, 9'sd172, 13'sd2512}, {4'sd4, 13'sd-2613, 12'sd-1644}, {13'sd-2301, 12'sd-1867, 12'sd1800}},
{{13'sd-2386, 9'sd148, 11'sd-845}, {12'sd-1752, 10'sd406, 13'sd2656}, {13'sd-2361, 12'sd-1578, 13'sd-2460}},
{{12'sd-1309, 12'sd-1919, 12'sd-1730}, {13'sd-2512, 9'sd133, 8'sd-67}, {13'sd2802, 10'sd414, 7'sd53}},
{{13'sd2632, 11'sd1002, 5'sd-14}, {12'sd-1984, 11'sd-653, 13'sd-2432}, {13'sd-2333, 13'sd2249, 13'sd2548}},
{{12'sd-1549, 12'sd-1937, 13'sd-2305}, {13'sd-2603, 11'sd-645, 11'sd921}, {13'sd-2555, 11'sd-932, 13'sd-2097}},
{{14'sd-4830, 12'sd-1665, 13'sd-4049}, {11'sd581, 11'sd-982, 10'sd-483}, {13'sd2223, 10'sd338, 12'sd-1505}},
{{13'sd2608, 13'sd-2063, 13'sd2284}, {11'sd-727, 13'sd2555, 12'sd-1852}, {13'sd2125, 11'sd-747, 11'sd-621}},
{{13'sd-2075, 13'sd-2628, 12'sd-1669}, {8'sd-96, 10'sd288, 12'sd-1503}, {13'sd2070, 13'sd2317, 12'sd-1062}},
{{12'sd-1105, 13'sd-2356, 11'sd991}, {9'sd-212, 12'sd-1499, 11'sd1012}, {13'sd3176, 11'sd570, 11'sd-684}},
{{11'sd526, 12'sd1651, 11'sd884}, {12'sd1361, 8'sd73, 12'sd-1807}, {13'sd2376, 12'sd-1296, 12'sd-1495}},
{{11'sd-938, 11'sd-806, 12'sd-1178}, {13'sd-2491, 13'sd-2988, 12'sd-1230}, {9'sd-202, 12'sd-1974, 13'sd2388}},
{{11'sd-717, 8'sd-105, 12'sd1042}, {12'sd1658, 12'sd-1411, 13'sd-2545}, {12'sd1179, 9'sd165, 7'sd43}},
{{12'sd-1677, 12'sd1470, 13'sd2445}, {13'sd-2723, 9'sd179, 11'sd752}, {11'sd-773, 10'sd403, 12'sd-1993}},
{{11'sd992, 12'sd-1060, 12'sd1593}, {12'sd-1171, 13'sd2052, 13'sd2248}, {12'sd-1435, 10'sd431, 13'sd-2820}},
{{11'sd-960, 9'sd159, 10'sd344}, {13'sd-2442, 13'sd-2219, 13'sd2360}, {10'sd-372, 8'sd72, 12'sd1150}},
{{12'sd1684, 12'sd-1790, 13'sd-2701}, {13'sd-2234, 12'sd1731, 10'sd463}, {12'sd1383, 11'sd-716, 13'sd-2172}},
{{12'sd1125, 12'sd-1435, 12'sd-1041}, {12'sd-1498, 12'sd-1418, 11'sd817}, {13'sd2715, 12'sd-1224, 12'sd1815}},
{{12'sd-1490, 12'sd1108, 13'sd3708}, {12'sd1946, 13'sd3501, 12'sd-1511}, {12'sd-1481, 8'sd106, 11'sd-774}},
{{10'sd-266, 11'sd622, 9'sd180}, {12'sd1201, 10'sd427, 9'sd-197}, {8'sd124, 13'sd-2779, 12'sd1870}},
{{12'sd-1670, 13'sd-2114, 13'sd-2781}, {9'sd250, 11'sd-630, 12'sd1755}, {9'sd252, 13'sd2128, 11'sd873}},
{{12'sd1270, 12'sd1177, 10'sd-447}, {13'sd2440, 13'sd-2078, 11'sd-920}, {11'sd-602, 12'sd-1741, 10'sd258}},
{{11'sd626, 12'sd-1917, 11'sd-768}, {10'sd423, 13'sd-2127, 8'sd-104}, {13'sd2137, 12'sd1626, 10'sd-333}},
{{10'sd337, 13'sd-2157, 11'sd532}, {13'sd2832, 12'sd1143, 12'sd1497}, {12'sd-1969, 10'sd451, 13'sd-2943}},
{{12'sd1389, 12'sd-1173, 12'sd1225}, {12'sd-1060, 6'sd-16, 12'sd1532}, {13'sd-2164, 10'sd-427, 12'sd1931}},
{{11'sd663, 13'sd2313, 12'sd1232}, {10'sd384, 12'sd-1954, 12'sd-1029}, {12'sd1697, 10'sd-414, 12'sd-1550}},
{{12'sd1300, 11'sd763, 8'sd111}, {12'sd-2011, 11'sd858, 11'sd651}, {12'sd1104, 12'sd1805, 13'sd2108}},
{{13'sd3479, 12'sd1301, 11'sd-815}, {13'sd2440, 10'sd256, 12'sd1835}, {12'sd-1356, 13'sd2051, 13'sd-2378}},
{{13'sd-2189, 11'sd-630, 12'sd1606}, {13'sd3013, 13'sd2812, 13'sd-2336}, {8'sd85, 6'sd-21, 13'sd2460}},
{{11'sd523, 12'sd-1151, 13'sd2310}, {12'sd1802, 12'sd1287, 11'sd-617}, {12'sd-1428, 12'sd1401, 12'sd1077}},
{{9'sd177, 11'sd-527, 13'sd2631}, {10'sd-327, 12'sd1743, 13'sd2443}, {11'sd-877, 12'sd1518, 11'sd679}},
{{12'sd1422, 12'sd1801, 13'sd-2318}, {12'sd-1510, 12'sd-1936, 11'sd906}, {12'sd1866, 11'sd-1001, 11'sd-814}},
{{12'sd1981, 12'sd-1826, 13'sd2982}, {13'sd-2367, 13'sd2316, 12'sd-1506}, {12'sd-1464, 12'sd-1454, 11'sd-714}},
{{12'sd-1989, 12'sd1934, 12'sd1725}, {13'sd-2612, 13'sd-2646, 12'sd-1585}, {12'sd1563, 10'sd-433, 13'sd-2128}},
{{10'sd-431, 13'sd-2130, 11'sd-660}, {12'sd1933, 11'sd640, 12'sd1556}, {11'sd-783, 10'sd304, 12'sd1644}},
{{13'sd2546, 12'sd-1370, 12'sd1705}, {10'sd-503, 12'sd-1185, 11'sd-790}, {7'sd32, 12'sd1666, 13'sd2336}},
{{13'sd2683, 13'sd2240, 12'sd-2020}, {11'sd-561, 12'sd1242, 12'sd-1787}, {12'sd1984, 13'sd2106, 7'sd-43}},
{{13'sd-2581, 10'sd441, 12'sd-1042}, {6'sd26, 10'sd386, 12'sd1088}, {12'sd1345, 12'sd1761, 9'sd196}},
{{12'sd1126, 12'sd1350, 9'sd-175}, {3'sd2, 12'sd1827, 12'sd1458}, {13'sd2283, 10'sd-349, 12'sd1601}},
{{12'sd1409, 12'sd1233, 13'sd2316}, {12'sd1763, 11'sd642, 12'sd1620}, {12'sd1512, 7'sd-40, 12'sd1865}},
{{13'sd2591, 13'sd-2352, 13'sd2201}, {11'sd-969, 10'sd-344, 12'sd-1876}, {12'sd-1737, 12'sd1832, 12'sd-1371}},
{{13'sd-2436, 12'sd-1453, 10'sd269}, {10'sd311, 13'sd2580, 11'sd697}, {12'sd1918, 13'sd3826, 12'sd1392}},
{{11'sd-694, 13'sd-2102, 9'sd243}, {7'sd-45, 8'sd-106, 12'sd-1984}, {11'sd-513, 11'sd-933, 13'sd-2148}},
{{12'sd-2022, 7'sd41, 12'sd-1815}, {7'sd-32, 12'sd-1884, 12'sd-1451}, {12'sd-1057, 7'sd-39, 12'sd-1143}},
{{10'sd-451, 11'sd532, 13'sd-2885}, {13'sd-2489, 11'sd-897, 9'sd138}, {11'sd-619, 12'sd1904, 13'sd-2209}},
{{11'sd932, 13'sd-2491, 11'sd1015}, {12'sd1216, 11'sd992, 13'sd-2679}, {11'sd729, 13'sd-2393, 13'sd-2232}},
{{13'sd-2524, 10'sd275, 13'sd-2643}, {11'sd599, 11'sd517, 12'sd-1176}, {13'sd2077, 12'sd2014, 12'sd-1485}},
{{13'sd-2392, 12'sd1213, 12'sd1385}, {12'sd-1180, 12'sd1628, 13'sd2314}, {13'sd2087, 13'sd2576, 11'sd966}},
{{12'sd-1254, 13'sd2916, 13'sd2595}, {13'sd2440, 12'sd1433, 11'sd559}, {11'sd-957, 12'sd-1467, 11'sd-1001}},
{{12'sd-1255, 12'sd1747, 12'sd1449}, {13'sd2073, 13'sd2614, 10'sd-425}, {12'sd1983, 11'sd768, 11'sd598}},
{{13'sd2338, 12'sd-1048, 11'sd565}, {12'sd1336, 12'sd1751, 12'sd-1775}, {11'sd-744, 13'sd-2140, 13'sd-2302}},
{{12'sd-1657, 11'sd608, 10'sd-465}, {12'sd-2029, 13'sd-2516, 9'sd244}, {11'sd-998, 12'sd-1247, 13'sd2272}},
{{12'sd-1237, 12'sd-1199, 9'sd-136}, {12'sd1114, 13'sd2067, 12'sd-1121}, {8'sd-77, 12'sd-1546, 12'sd-1585}}},
{
{{12'sd-1335, 12'sd-1755, 12'sd-1527}, {10'sd-400, 11'sd554, 12'sd1887}, {12'sd-1081, 11'sd512, 13'sd-2323}},
{{12'sd-1920, 12'sd1602, 13'sd2780}, {10'sd-453, 9'sd150, 12'sd-1349}, {13'sd-2458, 13'sd2191, 5'sd-11}},
{{12'sd-1328, 12'sd1268, 12'sd-1942}, {11'sd-598, 10'sd-508, 12'sd1795}, {13'sd2758, 13'sd3342, 11'sd629}},
{{13'sd2464, 11'sd-688, 13'sd2333}, {12'sd1336, 13'sd2129, 11'sd849}, {13'sd2400, 12'sd-1671, 12'sd-1199}},
{{12'sd-2027, 12'sd-2046, 12'sd1082}, {12'sd1769, 13'sd2380, 12'sd1449}, {12'sd1911, 13'sd2386, 10'sd496}},
{{12'sd-1956, 13'sd2413, 11'sd-721}, {11'sd-582, 12'sd2002, 13'sd2194}, {12'sd-1351, 13'sd2333, 12'sd2024}},
{{11'sd-888, 12'sd1824, 12'sd-1226}, {12'sd-1328, 13'sd-2265, 12'sd1381}, {13'sd2131, 13'sd-2084, 11'sd609}},
{{11'sd780, 10'sd-475, 12'sd-2041}, {13'sd2701, 11'sd854, 12'sd1107}, {13'sd-2569, 12'sd1635, 12'sd1686}},
{{11'sd-595, 12'sd1511, 11'sd963}, {10'sd266, 12'sd1177, 12'sd1456}, {13'sd2455, 12'sd1978, 12'sd-1760}},
{{13'sd-2363, 11'sd813, 13'sd2280}, {11'sd689, 13'sd2553, 13'sd2098}, {13'sd-2994, 9'sd-164, 12'sd1152}},
{{14'sd4609, 12'sd1516, 11'sd-808}, {13'sd3344, 12'sd1628, 11'sd804}, {9'sd167, 8'sd-118, 11'sd651}},
{{12'sd1599, 11'sd-988, 10'sd435}, {12'sd-1100, 13'sd2462, 11'sd-547}, {13'sd-2585, 12'sd1133, 13'sd-2199}},
{{9'sd-221, 12'sd-1725, 13'sd2560}, {12'sd-1666, 12'sd1972, 11'sd517}, {13'sd-2371, 10'sd372, 13'sd2563}},
{{11'sd845, 10'sd-432, 9'sd-225}, {12'sd1709, 10'sd426, 11'sd668}, {13'sd-2114, 13'sd-2511, 12'sd1473}},
{{12'sd1043, 12'sd-1861, 11'sd714}, {12'sd-1789, 12'sd1338, 11'sd-538}, {11'sd-564, 13'sd-2328, 12'sd-1846}},
{{10'sd-303, 10'sd446, 13'sd2478}, {12'sd1123, 11'sd619, 11'sd708}, {13'sd-2771, 13'sd2182, 13'sd2173}},
{{12'sd-1077, 11'sd984, 10'sd-306}, {9'sd-242, 11'sd-525, 11'sd953}, {10'sd-426, 12'sd-1736, 13'sd-2684}},
{{13'sd-2803, 13'sd-3427, 8'sd-84}, {9'sd-161, 10'sd-446, 11'sd951}, {12'sd1852, 13'sd2989, 11'sd-871}},
{{13'sd2640, 11'sd-791, 9'sd-143}, {13'sd2499, 10'sd-325, 12'sd1312}, {11'sd-732, 13'sd-2618, 12'sd1654}},
{{11'sd-623, 13'sd-2206, 12'sd-1122}, {11'sd-651, 12'sd-1357, 11'sd-913}, {12'sd1147, 12'sd1901, 13'sd-2461}},
{{9'sd-194, 10'sd336, 13'sd2352}, {13'sd2250, 12'sd1249, 11'sd908}, {13'sd2827, 12'sd-1647, 12'sd-1757}},
{{13'sd-2652, 12'sd1252, 11'sd-638}, {12'sd-1030, 10'sd-300, 10'sd276}, {12'sd-1111, 12'sd-1078, 11'sd855}},
{{11'sd789, 12'sd1536, 11'sd-836}, {9'sd-186, 8'sd-78, 13'sd-2748}, {10'sd260, 11'sd793, 13'sd2184}},
{{10'sd421, 12'sd-1195, 13'sd-2601}, {11'sd-550, 9'sd247, 12'sd2047}, {12'sd1505, 12'sd-1089, 11'sd569}},
{{13'sd-2883, 11'sd-681, 13'sd2316}, {12'sd-1205, 12'sd1516, 13'sd2725}, {12'sd1210, 12'sd1594, 11'sd-535}},
{{11'sd517, 12'sd-1694, 10'sd282}, {9'sd-188, 12'sd1758, 13'sd2171}, {10'sd333, 10'sd371, 13'sd-2307}},
{{12'sd-1674, 13'sd2778, 13'sd2299}, {13'sd-2292, 13'sd2833, 12'sd1211}, {12'sd-1647, 11'sd-943, 12'sd-1480}},
{{12'sd1653, 13'sd2552, 12'sd-1616}, {8'sd-96, 8'sd-117, 11'sd585}, {11'sd980, 10'sd494, 12'sd-1976}},
{{12'sd1759, 12'sd-1616, 13'sd2472}, {11'sd594, 11'sd938, 12'sd2047}, {8'sd71, 12'sd1640, 12'sd1097}},
{{13'sd2870, 12'sd1642, 11'sd568}, {13'sd2699, 9'sd148, 9'sd-172}, {10'sd-490, 11'sd696, 12'sd1936}},
{{13'sd-2485, 11'sd-964, 10'sd446}, {6'sd-19, 12'sd1111, 13'sd-2237}, {12'sd-2042, 13'sd2260, 9'sd142}},
{{13'sd2608, 12'sd1938, 10'sd470}, {12'sd-1551, 13'sd2101, 11'sd933}, {11'sd-883, 12'sd1886, 10'sd455}},
{{12'sd-1762, 13'sd-2557, 11'sd930}, {10'sd-273, 12'sd1970, 13'sd2372}, {12'sd-1902, 12'sd1070, 8'sd-87}},
{{10'sd-446, 7'sd-60, 12'sd1917}, {5'sd15, 10'sd369, 13'sd-2454}, {13'sd-2057, 12'sd1314, 10'sd-320}},
{{10'sd-416, 13'sd-2446, 12'sd1684}, {13'sd2100, 13'sd-2370, 11'sd846}, {12'sd-1822, 11'sd-724, 11'sd-893}},
{{12'sd-1440, 12'sd-1427, 11'sd966}, {13'sd2920, 9'sd133, 10'sd335}, {11'sd-527, 9'sd252, 7'sd50}},
{{13'sd-2245, 13'sd-2488, 12'sd-1757}, {13'sd2662, 12'sd-1683, 11'sd-863}, {12'sd-1785, 6'sd-19, 12'sd-1816}},
{{13'sd2488, 11'sd644, 11'sd701}, {12'sd1983, 11'sd769, 13'sd-2424}, {10'sd-510, 11'sd-549, 10'sd429}},
{{13'sd2678, 12'sd-1538, 9'sd-159}, {12'sd-1563, 11'sd576, 11'sd-803}, {11'sd700, 13'sd-2513, 12'sd-1248}},
{{12'sd-1994, 13'sd-2469, 10'sd-446}, {13'sd2234, 11'sd845, 12'sd1792}, {13'sd2286, 11'sd804, 10'sd408}},
{{12'sd1927, 13'sd-2060, 13'sd2987}, {12'sd-2034, 13'sd2333, 12'sd-1316}, {11'sd729, 10'sd-355, 13'sd-2510}},
{{11'sd588, 12'sd1052, 12'sd1815}, {12'sd-2011, 11'sd805, 12'sd1501}, {12'sd-1880, 13'sd2194, 11'sd-638}},
{{13'sd2682, 10'sd-376, 9'sd216}, {12'sd-2022, 13'sd2515, 12'sd1135}, {13'sd2636, 12'sd-1940, 13'sd2368}},
{{10'sd382, 12'sd-1571, 13'sd2472}, {13'sd2633, 12'sd-2021, 12'sd-1950}, {12'sd1323, 11'sd-588, 12'sd-1633}},
{{10'sd-426, 11'sd-710, 11'sd812}, {12'sd-1414, 12'sd-1725, 13'sd-2472}, {11'sd-905, 10'sd-380, 12'sd1343}},
{{13'sd-2787, 13'sd-2072, 10'sd-341}, {12'sd-1478, 10'sd277, 12'sd-1596}, {12'sd-1991, 12'sd-1929, 12'sd1024}},
{{13'sd2376, 11'sd-641, 6'sd-24}, {12'sd-1164, 13'sd2380, 13'sd-2756}, {12'sd1661, 11'sd942, 12'sd1608}},
{{12'sd1579, 10'sd-449, 12'sd1604}, {12'sd1221, 12'sd-1609, 13'sd-2580}, {9'sd150, 10'sd-507, 12'sd-1050}},
{{11'sd757, 12'sd1482, 12'sd1234}, {11'sd670, 12'sd-1532, 12'sd1451}, {11'sd-834, 11'sd748, 12'sd1477}},
{{13'sd2406, 13'sd-2158, 12'sd1402}, {13'sd2065, 8'sd120, 10'sd-409}, {10'sd-363, 13'sd-2758, 8'sd98}},
{{7'sd-60, 12'sd1319, 11'sd-1011}, {10'sd-511, 10'sd420, 13'sd2180}, {11'sd783, 12'sd-1828, 12'sd-1196}},
{{13'sd-2554, 13'sd2497, 12'sd1723}, {13'sd-2505, 13'sd-2341, 12'sd1172}, {9'sd177, 11'sd-727, 13'sd2422}},
{{12'sd-1394, 10'sd409, 13'sd-2931}, {11'sd-589, 5'sd-15, 13'sd-2264}, {12'sd1943, 13'sd2469, 11'sd-705}},
{{12'sd-1312, 12'sd-1754, 13'sd2216}, {12'sd-1127, 12'sd-1719, 11'sd545}, {12'sd1530, 11'sd607, 13'sd-2519}},
{{10'sd-269, 10'sd-354, 11'sd911}, {13'sd-2318, 12'sd1304, 12'sd-1400}, {13'sd-2584, 12'sd1788, 12'sd2032}},
{{12'sd-1285, 13'sd-2756, 12'sd1850}, {12'sd1308, 12'sd-1583, 12'sd-1385}, {12'sd-1971, 12'sd1485, 13'sd-2368}},
{{10'sd-314, 13'sd2457, 8'sd-70}, {11'sd-791, 11'sd-1005, 12'sd-1802}, {13'sd2328, 13'sd-2522, 13'sd2192}},
{{12'sd1130, 9'sd-150, 11'sd-1015}, {12'sd1895, 13'sd-2935, 12'sd-1642}, {13'sd2547, 11'sd852, 11'sd-555}},
{{12'sd1550, 11'sd722, 12'sd1073}, {11'sd973, 12'sd1943, 11'sd843}, {13'sd-2413, 12'sd-1060, 13'sd2583}},
{{13'sd-2316, 13'sd3016, 11'sd718}, {10'sd494, 9'sd167, 11'sd685}, {13'sd-2083, 12'sd1343, 13'sd2644}},
{{10'sd-388, 11'sd-835, 10'sd-510}, {13'sd2059, 7'sd-39, 11'sd872}, {12'sd1684, 12'sd1448, 11'sd-809}},
{{12'sd1141, 12'sd-1499, 9'sd129}, {7'sd39, 12'sd1874, 13'sd-2340}, {12'sd1836, 13'sd2121, 12'sd-1498}},
{{11'sd-897, 10'sd-373, 12'sd1065}, {13'sd-2950, 10'sd262, 12'sd1236}, {12'sd-1652, 10'sd-413, 13'sd-2922}},
{{13'sd-2961, 12'sd-1189, 13'sd-3272}, {13'sd-3106, 12'sd2031, 13'sd2099}, {11'sd524, 13'sd-2704, 13'sd2328}}},
{
{{12'sd-1360, 12'sd-1848, 12'sd-1526}, {12'sd1560, 10'sd485, 13'sd-2176}, {12'sd-1428, 11'sd-849, 11'sd-607}},
{{12'sd-1467, 13'sd2734, 12'sd-2000}, {13'sd-2082, 13'sd-2566, 13'sd2238}, {12'sd-1036, 11'sd-846, 10'sd-393}},
{{13'sd2520, 7'sd-44, 12'sd-1522}, {11'sd601, 10'sd-492, 12'sd1270}, {13'sd2585, 11'sd-891, 9'sd-151}},
{{13'sd-2920, 13'sd-2786, 13'sd-2293}, {10'sd-463, 10'sd-383, 13'sd-2946}, {11'sd936, 12'sd1986, 12'sd1388}},
{{12'sd-2018, 11'sd776, 12'sd-1414}, {11'sd-837, 7'sd54, 12'sd-1244}, {13'sd-2293, 12'sd1890, 12'sd-1893}},
{{13'sd2379, 13'sd-2445, 12'sd1213}, {12'sd-1439, 12'sd1929, 13'sd-2521}, {13'sd2485, 12'sd1193, 10'sd299}},
{{11'sd732, 11'sd-715, 10'sd-330}, {11'sd642, 12'sd-1482, 12'sd-1279}, {13'sd-2607, 11'sd-522, 13'sd2215}},
{{13'sd-2309, 13'sd-2463, 12'sd-1374}, {12'sd2033, 13'sd-2524, 11'sd538}, {4'sd-4, 8'sd-85, 12'sd1047}},
{{13'sd-2892, 12'sd1758, 10'sd-498}, {13'sd2218, 11'sd-606, 11'sd545}, {11'sd-810, 12'sd1202, 12'sd-1549}},
{{11'sd-728, 12'sd1692, 13'sd-2657}, {12'sd-1137, 12'sd1765, 9'sd-231}, {11'sd864, 13'sd-2184, 13'sd-2280}},
{{13'sd-2578, 11'sd-899, 13'sd2902}, {10'sd330, 12'sd1850, 10'sd363}, {10'sd361, 12'sd1135, 13'sd2098}},
{{12'sd-1898, 13'sd2183, 12'sd-1240}, {13'sd-2891, 12'sd1889, 12'sd1803}, {11'sd633, 13'sd2162, 11'sd655}},
{{12'sd-1421, 11'sd873, 9'sd147}, {13'sd2578, 12'sd1253, 12'sd-1199}, {11'sd620, 12'sd-1233, 12'sd-1835}},
{{12'sd-1666, 10'sd-446, 12'sd1719}, {12'sd1135, 12'sd-1251, 11'sd-576}, {10'sd-318, 13'sd-2256, 12'sd-1085}},
{{8'sd-100, 11'sd808, 13'sd2309}, {11'sd-735, 12'sd-1334, 11'sd1019}, {12'sd-1786, 9'sd187, 12'sd1991}},
{{9'sd-168, 12'sd-1832, 13'sd2487}, {13'sd2698, 12'sd1218, 10'sd390}, {12'sd1920, 13'sd2248, 11'sd715}},
{{13'sd2429, 12'sd-1559, 13'sd2336}, {13'sd3199, 12'sd1168, 13'sd-2783}, {12'sd-1600, 12'sd-1384, 12'sd-1210}},
{{13'sd2779, 11'sd-622, 11'sd526}, {13'sd2184, 11'sd808, 12'sd-1800}, {10'sd499, 13'sd-2792, 13'sd-3986}},
{{12'sd1076, 11'sd-832, 12'sd-1386}, {12'sd-1372, 13'sd-2735, 11'sd967}, {12'sd1054, 13'sd-2868, 13'sd2163}},
{{8'sd-93, 11'sd-892, 13'sd-2173}, {12'sd1082, 12'sd-1131, 13'sd-2553}, {10'sd450, 12'sd-1928, 12'sd1951}},
{{12'sd1731, 12'sd1951, 10'sd-447}, {13'sd2085, 12'sd1825, 11'sd641}, {11'sd1005, 12'sd-1140, 13'sd2891}},
{{13'sd2629, 11'sd-561, 12'sd1257}, {11'sd902, 12'sd-1803, 13'sd2967}, {11'sd-999, 11'sd-856, 13'sd3008}},
{{13'sd2304, 11'sd-613, 11'sd-627}, {11'sd769, 11'sd-665, 11'sd531}, {13'sd2537, 12'sd1867, 12'sd2008}},
{{12'sd1667, 12'sd-1537, 11'sd-634}, {13'sd-2658, 11'sd721, 10'sd-439}, {11'sd-766, 13'sd2719, 13'sd2338}},
{{13'sd2609, 10'sd455, 13'sd-2376}, {13'sd2408, 12'sd-1652, 10'sd-298}, {13'sd2227, 13'sd-2600, 12'sd-1732}},
{{13'sd-2839, 9'sd249, 12'sd-1750}, {11'sd721, 12'sd-1868, 12'sd-1667}, {8'sd81, 12'sd1178, 12'sd1648}},
{{12'sd-1176, 13'sd-2402, 11'sd-596}, {11'sd-512, 13'sd-2452, 12'sd1040}, {13'sd-2699, 12'sd1508, 13'sd-2493}},
{{10'sd-384, 12'sd-1629, 11'sd601}, {9'sd181, 13'sd-2687, 12'sd-1773}, {12'sd-1862, 11'sd819, 13'sd-2812}},
{{13'sd2615, 10'sd461, 12'sd1847}, {10'sd-374, 9'sd193, 13'sd-2209}, {12'sd-1200, 13'sd-2606, 10'sd347}},
{{12'sd-1808, 11'sd795, 13'sd-2451}, {12'sd1113, 11'sd974, 11'sd754}, {12'sd1587, 13'sd2276, 11'sd727}},
{{12'sd1858, 12'sd1957, 11'sd708}, {12'sd-1302, 13'sd2317, 11'sd576}, {12'sd-1498, 13'sd2812, 10'sd-447}},
{{12'sd-1663, 12'sd-2009, 12'sd-1037}, {12'sd1820, 13'sd-2567, 12'sd-1081}, {12'sd-2031, 10'sd-413, 12'sd-1328}},
{{8'sd-96, 13'sd2292, 12'sd-1132}, {13'sd2663, 9'sd199, 13'sd2468}, {10'sd476, 11'sd-630, 10'sd400}},
{{12'sd-1234, 10'sd-384, 13'sd-2241}, {12'sd-1326, 12'sd1089, 9'sd218}, {13'sd2574, 9'sd-189, 12'sd-1072}},
{{12'sd-1516, 13'sd-2104, 11'sd-591}, {12'sd-1099, 12'sd-1516, 13'sd2107}, {10'sd-374, 12'sd1126, 12'sd-1681}},
{{12'sd1770, 12'sd-1692, 13'sd-2458}, {11'sd585, 13'sd-2772, 10'sd-317}, {9'sd255, 12'sd1901, 12'sd-1857}},
{{12'sd-1619, 11'sd935, 12'sd1659}, {13'sd2130, 10'sd-381, 13'sd2254}, {12'sd-1439, 13'sd-2143, 12'sd1555}},
{{13'sd2269, 13'sd-2254, 12'sd1424}, {10'sd-397, 9'sd-187, 12'sd-2045}, {11'sd-955, 13'sd-2368, 12'sd-1282}},
{{12'sd-1455, 11'sd-612, 6'sd-28}, {10'sd500, 10'sd-294, 11'sd-970}, {13'sd-2068, 12'sd1814, 13'sd-2288}},
{{10'sd-388, 12'sd1630, 8'sd-79}, {11'sd-905, 9'sd-180, 11'sd-626}, {13'sd-2455, 11'sd610, 13'sd2406}},
{{11'sd-912, 10'sd-489, 9'sd-159}, {12'sd1224, 13'sd3155, 11'sd-927}, {10'sd376, 12'sd1667, 13'sd-2815}},
{{13'sd2378, 11'sd829, 11'sd551}, {12'sd1177, 12'sd-1628, 8'sd-120}, {12'sd-1226, 9'sd215, 10'sd-393}},
{{10'sd352, 9'sd-250, 10'sd-407}, {12'sd-1770, 13'sd2156, 13'sd-2295}, {12'sd-2006, 11'sd-687, 11'sd751}},
{{13'sd-2544, 12'sd1746, 12'sd1506}, {10'sd324, 9'sd-172, 12'sd-1662}, {12'sd1073, 12'sd1336, 6'sd-17}},
{{10'sd-383, 11'sd-885, 10'sd-310}, {13'sd2552, 13'sd2438, 10'sd-269}, {8'sd127, 12'sd1063, 10'sd-480}},
{{11'sd-826, 10'sd-373, 12'sd1932}, {9'sd-253, 12'sd1057, 13'sd2240}, {13'sd2666, 13'sd-2279, 12'sd-1678}},
{{13'sd2507, 12'sd-1603, 13'sd3046}, {12'sd-1919, 11'sd932, 13'sd2169}, {13'sd2079, 9'sd155, 13'sd-2099}},
{{13'sd-2617, 12'sd1789, 12'sd1388}, {12'sd-1346, 11'sd800, 11'sd1017}, {11'sd928, 13'sd-2304, 10'sd-334}},
{{13'sd2456, 12'sd-1848, 12'sd-1081}, {11'sd597, 10'sd395, 12'sd-1662}, {11'sd-793, 13'sd-2364, 13'sd-2211}},
{{13'sd-2673, 10'sd303, 11'sd-921}, {12'sd1680, 12'sd1965, 13'sd2156}, {13'sd2259, 13'sd2498, 13'sd2338}},
{{12'sd-1913, 12'sd1586, 12'sd-1069}, {12'sd1544, 12'sd-1243, 10'sd484}, {13'sd-2357, 12'sd1093, 12'sd1875}},
{{11'sd1014, 11'sd-514, 7'sd-47}, {9'sd182, 9'sd-163, 12'sd-1848}, {12'sd-1048, 12'sd2030, 10'sd-391}},
{{11'sd-747, 13'sd2337, 13'sd3057}, {12'sd2032, 12'sd1960, 11'sd-914}, {12'sd-1151, 13'sd-2996, 12'sd-1547}},
{{9'sd-132, 13'sd3034, 12'sd-1803}, {11'sd735, 12'sd-1210, 7'sd59}, {11'sd944, 11'sd-734, 13'sd-2441}},
{{11'sd789, 12'sd1822, 12'sd-1698}, {11'sd-888, 12'sd-1623, 9'sd-208}, {12'sd1478, 13'sd2178, 13'sd3051}},
{{10'sd434, 12'sd-1074, 9'sd177}, {11'sd-951, 12'sd1230, 13'sd2445}, {10'sd402, 7'sd35, 13'sd2754}},
{{12'sd-1979, 11'sd-656, 10'sd298}, {10'sd-393, 12'sd-1769, 12'sd1276}, {13'sd-2373, 11'sd-924, 12'sd2003}},
{{13'sd2236, 13'sd2192, 10'sd-325}, {11'sd650, 12'sd1202, 13'sd2114}, {12'sd-1155, 12'sd-1159, 11'sd-625}},
{{10'sd434, 12'sd1121, 12'sd1398}, {12'sd-1796, 10'sd303, 9'sd-213}, {8'sd-104, 11'sd1018, 10'sd311}},
{{12'sd1919, 12'sd-1117, 12'sd-1740}, {11'sd-537, 11'sd-985, 12'sd-1429}, {12'sd1653, 12'sd1350, 13'sd-2406}},
{{11'sd901, 11'sd768, 12'sd-1903}, {12'sd-1354, 12'sd1730, 9'sd170}, {13'sd2607, 11'sd976, 12'sd1512}},
{{12'sd-1915, 12'sd1950, 13'sd-2258}, {10'sd436, 12'sd-1068, 12'sd1776}, {13'sd2166, 12'sd1537, 11'sd-740}},
{{12'sd-1215, 11'sd-692, 11'sd906}, {13'sd-2306, 13'sd-2255, 12'sd1137}, {11'sd-614, 12'sd-1466, 13'sd2221}},
{{8'sd-64, 10'sd-482, 13'sd2308}, {12'sd1385, 11'sd551, 11'sd-929}, {12'sd-1652, 13'sd-2762, 12'sd-1542}}},
{
{{12'sd1651, 11'sd-533, 11'sd910}, {9'sd220, 12'sd2013, 13'sd3050}, {12'sd-1099, 9'sd-143, 10'sd432}},
{{11'sd-924, 11'sd-638, 11'sd571}, {12'sd-1541, 12'sd-2037, 9'sd239}, {11'sd-742, 11'sd-564, 13'sd-2782}},
{{11'sd763, 7'sd63, 10'sd-386}, {12'sd-1404, 13'sd-2469, 10'sd-466}, {13'sd-3006, 12'sd1308, 12'sd1831}},
{{11'sd-903, 12'sd1915, 13'sd-2539}, {12'sd1554, 12'sd-1180, 12'sd-1130}, {12'sd1408, 7'sd-59, 12'sd-1546}},
{{12'sd1784, 13'sd-2815, 12'sd1148}, {13'sd-2407, 11'sd-730, 11'sd650}, {12'sd-1142, 7'sd63, 6'sd-20}},
{{12'sd-1485, 13'sd-2321, 12'sd1792}, {13'sd-2455, 10'sd-504, 12'sd-1207}, {12'sd-1130, 12'sd-1036, 13'sd-2670}},
{{13'sd3622, 11'sd848, 11'sd998}, {11'sd918, 13'sd2887, 11'sd571}, {12'sd1149, 13'sd2886, 8'sd111}},
{{12'sd1365, 13'sd-2864, 13'sd2715}, {10'sd307, 13'sd-3593, 11'sd585}, {12'sd-1484, 11'sd-968, 13'sd-2867}},
{{11'sd-856, 12'sd-1258, 12'sd-1243}, {10'sd-264, 8'sd-119, 13'sd-2916}, {12'sd-1467, 9'sd-206, 12'sd-1593}},
{{11'sd-933, 11'sd969, 13'sd-2359}, {13'sd2921, 9'sd-158, 13'sd-2372}, {12'sd-1976, 12'sd1165, 10'sd-501}},
{{14'sd4863, 10'sd347, 11'sd624}, {13'sd3766, 13'sd3447, 12'sd-1806}, {12'sd-1701, 11'sd993, 13'sd-3721}},
{{12'sd-1882, 6'sd20, 9'sd-247}, {13'sd-2356, 13'sd-2641, 13'sd-2271}, {12'sd1442, 13'sd-3861, 12'sd1377}},
{{14'sd4559, 11'sd659, 13'sd2289}, {12'sd-1300, 11'sd987, 13'sd2052}, {10'sd267, 12'sd-1915, 14'sd4667}},
{{12'sd-1125, 10'sd365, 12'sd1116}, {13'sd-2076, 13'sd2433, 12'sd-1228}, {11'sd-894, 13'sd-2473, 13'sd-2821}},
{{12'sd-1326, 13'sd-2354, 12'sd1081}, {12'sd1619, 9'sd248, 11'sd-572}, {13'sd2659, 12'sd1533, 13'sd-2669}},
{{13'sd2280, 11'sd747, 13'sd2280}, {12'sd1559, 10'sd439, 13'sd2108}, {13'sd2761, 11'sd750, 11'sd570}},
{{13'sd2092, 11'sd-785, 13'sd2811}, {12'sd-1798, 12'sd-1535, 13'sd2780}, {9'sd214, 7'sd53, 12'sd1638}},
{{6'sd26, 12'sd-1109, 11'sd-713}, {13'sd-3084, 11'sd-794, 12'sd-1548}, {13'sd-2908, 13'sd-2089, 10'sd268}},
{{12'sd-1157, 13'sd2233, 11'sd-660}, {13'sd-2287, 13'sd2357, 12'sd-1271}, {7'sd-47, 13'sd-2201, 11'sd967}},
{{12'sd-1776, 11'sd-735, 12'sd-1582}, {13'sd-2576, 13'sd3084, 13'sd-2292}, {8'sd78, 7'sd40, 11'sd921}},
{{12'sd2020, 9'sd-240, 13'sd-2272}, {12'sd-1528, 11'sd-781, 12'sd-1890}, {13'sd2378, 13'sd2049, 11'sd-733}},
{{8'sd-122, 11'sd-516, 12'sd1525}, {12'sd-1027, 13'sd3077, 12'sd-1351}, {7'sd56, 12'sd1660, 13'sd-2511}},
{{12'sd-1678, 10'sd-437, 12'sd1323}, {10'sd306, 13'sd-2271, 13'sd2111}, {13'sd2447, 12'sd-1979, 12'sd-1221}},
{{13'sd2301, 10'sd288, 11'sd-849}, {12'sd-1506, 12'sd1906, 11'sd1003}, {13'sd2842, 11'sd-792, 8'sd-118}},
{{12'sd-1818, 13'sd-2398, 12'sd-1548}, {13'sd2093, 13'sd-3681, 10'sd-465}, {13'sd-2877, 12'sd-1235, 12'sd1516}},
{{12'sd-1948, 11'sd694, 12'sd-1680}, {12'sd2019, 12'sd-1740, 13'sd2674}, {12'sd-1320, 13'sd2465, 11'sd576}},
{{13'sd2076, 13'sd2242, 13'sd-2119}, {13'sd-2719, 13'sd2694, 13'sd-2487}, {12'sd-1191, 13'sd2157, 13'sd-3521}},
{{11'sd963, 12'sd1659, 11'sd946}, {13'sd2475, 12'sd-1760, 13'sd-2118}, {12'sd-1206, 13'sd-2330, 9'sd-242}},
{{12'sd1963, 13'sd2873, 12'sd-2025}, {12'sd1302, 13'sd2505, 13'sd-2088}, {12'sd-1963, 13'sd2864, 11'sd752}},
{{12'sd1463, 12'sd-1717, 12'sd-1718}, {13'sd2369, 11'sd646, 12'sd1634}, {13'sd3005, 11'sd834, 12'sd1038}},
{{13'sd2063, 3'sd-2, 11'sd550}, {12'sd1650, 13'sd2388, 11'sd888}, {9'sd231, 13'sd2675, 13'sd2582}},
{{7'sd62, 13'sd-2812, 12'sd1101}, {12'sd1288, 12'sd-1327, 11'sd-681}, {13'sd-2291, 13'sd-2815, 11'sd-805}},
{{13'sd2119, 12'sd1744, 13'sd3047}, {13'sd2834, 11'sd516, 11'sd-632}, {11'sd910, 12'sd2033, 11'sd-992}},
{{10'sd-354, 13'sd-2614, 12'sd-1549}, {11'sd-837, 12'sd-1229, 12'sd1807}, {11'sd-1023, 13'sd2358, 10'sd316}},
{{12'sd-1898, 13'sd2448, 10'sd356}, {12'sd1350, 13'sd2406, 13'sd-2493}, {12'sd-1797, 10'sd410, 11'sd832}},
{{12'sd-1391, 9'sd-167, 11'sd559}, {12'sd1070, 11'sd-795, 12'sd-1681}, {10'sd-439, 10'sd-421, 12'sd-1746}},
{{12'sd-1057, 13'sd-2078, 10'sd-498}, {12'sd-1919, 13'sd-2680, 12'sd-1971}, {9'sd-214, 11'sd826, 13'sd-2468}},
{{13'sd-3226, 10'sd399, 13'sd2873}, {13'sd2424, 10'sd449, 10'sd257}, {13'sd-3784, 9'sd236, 13'sd-2163}},
{{11'sd-864, 13'sd3151, 11'sd852}, {13'sd2376, 9'sd206, 8'sd120}, {12'sd-1169, 13'sd-2914, 12'sd-1511}},
{{10'sd-277, 13'sd3448, 13'sd2671}, {13'sd2248, 10'sd-392, 11'sd767}, {10'sd-413, 13'sd-2679, 12'sd1495}},
{{13'sd2187, 10'sd356, 13'sd2135}, {12'sd-1272, 11'sd837, 12'sd1070}, {9'sd190, 10'sd-380, 12'sd-1359}},
{{13'sd2288, 10'sd289, 12'sd1486}, {11'sd-646, 12'sd-1535, 12'sd1950}, {11'sd540, 13'sd-3304, 12'sd1731}},
{{12'sd-1435, 12'sd-1809, 12'sd2005}, {10'sd383, 12'sd-2043, 13'sd-2719}, {13'sd-2095, 12'sd2015, 6'sd21}},
{{12'sd-1870, 13'sd2180, 9'sd-163}, {12'sd-1785, 12'sd1550, 11'sd1013}, {12'sd1354, 11'sd873, 12'sd1234}},
{{13'sd-2803, 8'sd-108, 13'sd-2538}, {12'sd1725, 12'sd1501, 13'sd-2977}, {12'sd-1075, 12'sd1305, 12'sd-1064}},
{{12'sd1342, 11'sd-862, 11'sd-829}, {13'sd2527, 12'sd1658, 12'sd1328}, {12'sd-1442, 12'sd-1642, 11'sd803}},
{{13'sd2860, 13'sd-2140, 10'sd440}, {9'sd251, 13'sd2595, 12'sd1595}, {7'sd45, 13'sd3047, 13'sd2955}},
{{12'sd-1141, 12'sd-2040, 12'sd-1498}, {11'sd966, 9'sd223, 12'sd-1276}, {11'sd-814, 11'sd-735, 10'sd286}},
{{7'sd49, 12'sd-1072, 13'sd2131}, {13'sd-2131, 10'sd-279, 13'sd2280}, {10'sd-256, 12'sd1846, 7'sd63}},
{{11'sd-849, 13'sd3178, 12'sd-1630}, {11'sd-540, 7'sd33, 12'sd-1317}, {13'sd2691, 9'sd195, 13'sd-2410}},
{{13'sd-2405, 10'sd450, 9'sd181}, {10'sd307, 12'sd1218, 12'sd1424}, {12'sd2016, 9'sd227, 11'sd-573}},
{{13'sd2871, 11'sd-742, 12'sd1235}, {13'sd-2381, 12'sd1274, 12'sd-1522}, {11'sd-695, 13'sd2742, 12'sd-1151}},
{{13'sd-2200, 11'sd588, 6'sd25}, {10'sd-438, 13'sd-2774, 13'sd-2626}, {13'sd-2844, 12'sd-1662, 14'sd-4667}},
{{11'sd-617, 12'sd1864, 11'sd-987}, {12'sd1587, 12'sd-1740, 12'sd1798}, {11'sd-767, 10'sd-385, 13'sd2068}},
{{10'sd441, 12'sd1209, 9'sd-193}, {9'sd-237, 12'sd-1583, 13'sd2655}, {9'sd151, 12'sd1603, 13'sd2389}},
{{12'sd-1542, 12'sd-2032, 12'sd-1127}, {12'sd-1165, 11'sd-975, 12'sd-1056}, {12'sd1271, 13'sd2481, 12'sd-1716}},
{{8'sd-119, 12'sd-1638, 12'sd-1763}, {11'sd961, 12'sd-1537, 13'sd-2480}, {9'sd236, 8'sd-95, 13'sd2664}},
{{13'sd3635, 12'sd-1226, 13'sd2449}, {9'sd230, 12'sd-1239, 10'sd-397}, {13'sd-3690, 12'sd-1701, 11'sd-537}},
{{12'sd1776, 11'sd534, 12'sd1825}, {12'sd-1899, 10'sd-369, 13'sd-2408}, {13'sd3488, 14'sd4419, 12'sd1265}},
{{12'sd1944, 12'sd1590, 13'sd2357}, {13'sd2134, 12'sd1600, 13'sd-2563}, {13'sd-2525, 12'sd-1193, 11'sd684}},
{{12'sd1181, 13'sd-2191, 9'sd209}, {9'sd165, 13'sd-2993, 12'sd-1318}, {12'sd1774, 12'sd1753, 11'sd-921}},
{{11'sd-916, 12'sd1547, 11'sd994}, {13'sd-2404, 12'sd1162, 13'sd2107}, {13'sd2498, 13'sd2404, 13'sd-2349}},
{{11'sd-801, 12'sd-1669, 13'sd-2351}, {13'sd-2150, 12'sd-1915, 10'sd463}, {12'sd-1891, 11'sd562, 12'sd-1557}},
{{9'sd204, 13'sd-2062, 13'sd2366}, {11'sd-795, 12'sd1191, 11'sd655}, {12'sd1309, 12'sd1471, 13'sd2982}}},
{
{{11'sd763, 12'sd-1973, 13'sd-2361}, {9'sd-203, 13'sd-2781, 13'sd2316}, {12'sd-1984, 5'sd-9, 12'sd1717}},
{{13'sd-2610, 11'sd612, 8'sd-76}, {12'sd2013, 7'sd-40, 11'sd-944}, {10'sd-455, 8'sd-95, 13'sd-2677}},
{{6'sd27, 12'sd-1588, 12'sd-1732}, {12'sd-1377, 8'sd109, 13'sd3579}, {13'sd3179, 12'sd-1629, 13'sd2608}},
{{11'sd-667, 12'sd1382, 12'sd1343}, {12'sd-1465, 9'sd-177, 9'sd240}, {11'sd646, 10'sd-484, 9'sd168}},
{{7'sd43, 12'sd1257, 11'sd-557}, {12'sd-1245, 13'sd2369, 10'sd505}, {7'sd61, 10'sd-503, 10'sd-391}},
{{13'sd2704, 12'sd-1194, 8'sd-125}, {13'sd2074, 13'sd-2367, 13'sd2873}, {13'sd2973, 10'sd270, 11'sd823}},
{{12'sd1133, 9'sd154, 12'sd1772}, {9'sd179, 13'sd-2065, 12'sd-1538}, {13'sd2127, 13'sd2658, 11'sd-589}},
{{13'sd-2324, 13'sd-2228, 10'sd274}, {8'sd122, 13'sd-3154, 11'sd938}, {13'sd2399, 12'sd-1833, 13'sd2251}},
{{12'sd-1514, 13'sd-2740, 11'sd613}, {12'sd-1536, 12'sd-1550, 11'sd903}, {13'sd3288, 11'sd817, 13'sd2650}},
{{11'sd-974, 10'sd-369, 11'sd617}, {11'sd636, 10'sd-428, 8'sd-94}, {12'sd-1286, 11'sd-994, 13'sd-2477}},
{{14'sd5661, 14'sd5316, 13'sd3808}, {10'sd-447, 13'sd2685, 11'sd1009}, {10'sd-425, 12'sd1657, 12'sd-1880}},
{{10'sd349, 10'sd281, 12'sd1573}, {10'sd-258, 12'sd1975, 11'sd754}, {12'sd-1967, 12'sd1544, 7'sd47}},
{{11'sd-655, 13'sd-3177, 12'sd-1647}, {13'sd-2429, 9'sd176, 11'sd965}, {12'sd-1652, 13'sd-2839, 12'sd-1415}},
{{13'sd2311, 11'sd512, 12'sd-1615}, {10'sd-300, 12'sd1772, 12'sd1234}, {13'sd-2614, 11'sd583, 8'sd-127}},
{{11'sd776, 12'sd-1186, 12'sd-1825}, {12'sd1835, 11'sd1011, 12'sd-1713}, {13'sd-2604, 9'sd-181, 9'sd174}},
{{12'sd-1385, 11'sd922, 11'sd-759}, {10'sd325, 13'sd-2582, 9'sd-207}, {10'sd274, 12'sd1289, 11'sd-1011}},
{{13'sd-2190, 13'sd-2211, 11'sd-1017}, {10'sd-289, 13'sd-3279, 9'sd-167}, {12'sd-1855, 12'sd1082, 11'sd-594}},
{{13'sd-3324, 13'sd-2638, 11'sd-644}, {12'sd1882, 12'sd-1127, 13'sd-3106}, {11'sd851, 13'sd3212, 12'sd-1407}},
{{11'sd-564, 13'sd2086, 9'sd237}, {13'sd-2622, 13'sd-2052, 12'sd1963}, {6'sd-30, 12'sd-1362, 13'sd-2537}},
{{13'sd2533, 9'sd199, 8'sd91}, {13'sd2731, 10'sd-267, 13'sd-3423}, {12'sd1746, 11'sd-950, 13'sd-2208}},
{{13'sd-2664, 11'sd-907, 11'sd531}, {12'sd-1755, 12'sd-1951, 11'sd-687}, {11'sd612, 9'sd-220, 11'sd-531}},
{{13'sd-2403, 11'sd1022, 13'sd3647}, {13'sd-2059, 10'sd-477, 13'sd2096}, {12'sd1406, 11'sd-611, 7'sd44}},
{{12'sd-1199, 10'sd317, 12'sd1827}, {11'sd-784, 12'sd-2003, 10'sd431}, {12'sd1609, 12'sd-1731, 12'sd-1706}},
{{11'sd-1004, 10'sd280, 11'sd-544}, {13'sd2465, 12'sd1406, 9'sd-128}, {8'sd-93, 8'sd95, 12'sd1321}},
{{4'sd-5, 13'sd-2890, 13'sd2848}, {13'sd-2192, 10'sd-421, 5'sd-11}, {14'sd4304, 12'sd1997, 14'sd4412}},
{{13'sd2678, 13'sd-2185, 12'sd-1197}, {12'sd1732, 12'sd-1060, 9'sd-187}, {12'sd1678, 12'sd-1766, 13'sd-2414}},
{{11'sd934, 13'sd-2053, 11'sd960}, {11'sd1005, 8'sd-100, 11'sd971}, {12'sd1865, 12'sd1768, 13'sd-2513}},
{{11'sd821, 12'sd-1108, 13'sd-2306}, {11'sd-633, 12'sd1198, 12'sd-1171}, {10'sd355, 9'sd-255, 12'sd-1329}},
{{11'sd513, 13'sd3071, 13'sd-2117}, {12'sd-1184, 10'sd345, 12'sd1601}, {12'sd1599, 11'sd-846, 13'sd-2949}},
{{11'sd-974, 11'sd-841, 12'sd1656}, {11'sd-888, 13'sd2131, 10'sd378}, {12'sd-1959, 13'sd-2655, 10'sd-415}},
{{12'sd-1263, 8'sd65, 11'sd-518}, {12'sd-1570, 10'sd388, 11'sd882}, {12'sd-1201, 12'sd-1376, 9'sd154}},
{{11'sd-569, 13'sd-3344, 13'sd-3328}, {12'sd1216, 13'sd-3006, 13'sd-2173}, {11'sd944, 11'sd-793, 8'sd-79}},
{{11'sd972, 12'sd-2046, 11'sd-641}, {12'sd1411, 8'sd107, 12'sd1757}, {11'sd-558, 12'sd1731, 12'sd1259}},
{{12'sd-1213, 12'sd1278, 12'sd1431}, {11'sd888, 11'sd-532, 13'sd2749}, {10'sd311, 13'sd2150, 9'sd-187}},
{{12'sd2030, 10'sd379, 12'sd-1176}, {11'sd539, 13'sd2364, 10'sd313}, {12'sd-1157, 10'sd468, 11'sd915}},
{{11'sd-986, 12'sd-1372, 10'sd295}, {9'sd-237, 13'sd-2487, 12'sd-1660}, {11'sd-1002, 13'sd2432, 10'sd-507}},
{{10'sd501, 13'sd2231, 12'sd1618}, {12'sd1062, 12'sd-2026, 12'sd-1203}, {12'sd1843, 11'sd-746, 12'sd-1528}},
{{10'sd-504, 12'sd1187, 12'sd-1171}, {4'sd-6, 13'sd2373, 13'sd-2108}, {11'sd-943, 12'sd-1414, 12'sd1203}},
{{13'sd2952, 10'sd-331, 13'sd2108}, {13'sd2331, 13'sd-3162, 13'sd-2649}, {13'sd2227, 13'sd-2506, 11'sd-672}},
{{12'sd-1427, 12'sd1911, 11'sd-784}, {12'sd-1220, 13'sd2344, 12'sd1682}, {12'sd1369, 11'sd566, 12'sd1653}},
{{12'sd-1048, 12'sd1476, 12'sd-1365}, {13'sd2571, 13'sd2824, 10'sd429}, {12'sd1880, 12'sd-2026, 11'sd-550}},
{{13'sd-2375, 10'sd485, 13'sd-2343}, {11'sd762, 11'sd515, 10'sd355}, {12'sd-1804, 10'sd-409, 11'sd-851}},
{{12'sd-1451, 13'sd2097, 12'sd1057}, {12'sd-1922, 13'sd2580, 12'sd1849}, {7'sd-45, 10'sd-305, 12'sd-1654}},
{{11'sd861, 6'sd23, 11'sd836}, {11'sd941, 11'sd-769, 13'sd2436}, {12'sd1357, 11'sd-853, 11'sd518}},
{{11'sd530, 7'sd-45, 13'sd2325}, {12'sd1514, 11'sd-834, 11'sd-764}, {11'sd545, 11'sd867, 11'sd843}},
{{12'sd1513, 11'sd792, 13'sd2476}, {13'sd3111, 12'sd1052, 12'sd-1901}, {12'sd-1807, 10'sd310, 13'sd-2085}},
{{10'sd463, 13'sd2478, 12'sd-1854}, {13'sd-2919, 12'sd-1237, 11'sd589}, {10'sd-283, 12'sd1121, 12'sd-1222}},
{{12'sd-1465, 12'sd1787, 12'sd-1215}, {9'sd220, 12'sd-1241, 10'sd-378}, {12'sd-1779, 13'sd2530, 12'sd-1297}},
{{13'sd-2265, 11'sd-876, 10'sd411}, {10'sd383, 12'sd1252, 9'sd-201}, {11'sd-700, 11'sd549, 12'sd1605}},
{{10'sd-272, 13'sd2460, 11'sd661}, {8'sd110, 13'sd-2968, 13'sd-2349}, {13'sd2052, 13'sd-2896, 8'sd-116}},
{{12'sd-1753, 11'sd891, 12'sd1716}, {13'sd-2991, 13'sd-2167, 12'sd-1222}, {11'sd-971, 12'sd-1374, 12'sd-1068}},
{{12'sd-1060, 12'sd1355, 12'sd2030}, {10'sd395, 8'sd125, 13'sd-2276}, {12'sd-1188, 10'sd375, 12'sd1252}},
{{12'sd-1153, 13'sd2221, 12'sd-1064}, {10'sd-301, 12'sd1451, 13'sd-2089}, {10'sd-499, 12'sd1517, 12'sd1699}},
{{12'sd-2013, 12'sd1862, 13'sd-2488}, {12'sd1026, 12'sd1812, 12'sd-1551}, {11'sd998, 10'sd369, 8'sd127}},
{{12'sd1799, 10'sd-339, 11'sd-792}, {12'sd1312, 12'sd1990, 12'sd-1335}, {12'sd-1225, 13'sd-2334, 13'sd-2201}},
{{12'sd1822, 11'sd-670, 12'sd-1245}, {12'sd1445, 12'sd-1922, 12'sd1532}, {11'sd987, 11'sd-606, 13'sd2150}},
{{12'sd1096, 11'sd-778, 12'sd-1561}, {12'sd-1456, 12'sd-1370, 10'sd438}, {8'sd-75, 10'sd-290, 13'sd2628}},
{{13'sd2298, 13'sd-2613, 12'sd1044}, {12'sd-1495, 13'sd-2605, 10'sd-327}, {13'sd3125, 12'sd1122, 13'sd3444}},
{{13'sd2180, 11'sd-676, 11'sd-518}, {11'sd-571, 13'sd3330, 10'sd-505}, {13'sd3122, 13'sd4003, 12'sd1225}},
{{12'sd1443, 11'sd-659, 11'sd845}, {13'sd-2309, 12'sd1498, 13'sd-2959}, {11'sd737, 6'sd-29, 11'sd-713}},
{{13'sd-3049, 12'sd-1192, 13'sd-2254}, {12'sd1046, 13'sd-2841, 12'sd1699}, {13'sd2495, 13'sd2234, 12'sd-1395}},
{{12'sd-1079, 12'sd1496, 11'sd750}, {12'sd1865, 12'sd1312, 12'sd-1526}, {13'sd-2751, 9'sd191, 11'sd948}},
{{13'sd2654, 10'sd-461, 13'sd-2288}, {5'sd10, 12'sd1532, 12'sd-1917}, {13'sd2533, 12'sd-1642, 11'sd-656}},
{{9'sd197, 10'sd262, 11'sd808}, {10'sd-334, 10'sd-511, 4'sd-6}, {8'sd-87, 12'sd1297, 13'sd2544}}},
{
{{10'sd399, 11'sd-715, 12'sd1400}, {12'sd-1207, 13'sd-2962, 12'sd-1639}, {10'sd381, 12'sd-1645, 12'sd-1294}},
{{13'sd-2227, 11'sd516, 13'sd2831}, {13'sd-2150, 11'sd852, 12'sd1393}, {12'sd-1652, 12'sd1473, 12'sd-1565}},
{{12'sd-1537, 11'sd585, 13'sd3077}, {13'sd-2084, 9'sd-151, 13'sd3964}, {11'sd-944, 11'sd947, 12'sd-1222}},
{{12'sd-1733, 13'sd2719, 12'sd1853}, {12'sd1390, 12'sd1046, 10'sd-414}, {11'sd-714, 10'sd382, 13'sd-2863}},
{{11'sd-604, 10'sd-360, 12'sd1367}, {13'sd-3186, 13'sd-2645, 12'sd-2001}, {12'sd-1299, 13'sd-2355, 12'sd1092}},
{{12'sd-1722, 13'sd2140, 11'sd976}, {12'sd-1591, 12'sd1910, 11'sd991}, {11'sd-521, 13'sd2621, 12'sd-1286}},
{{11'sd774, 12'sd-1632, 13'sd2170}, {8'sd-111, 12'sd-1890, 12'sd-1517}, {9'sd146, 11'sd-886, 13'sd2888}},
{{13'sd2760, 12'sd-1433, 12'sd-1291}, {12'sd1096, 12'sd1664, 13'sd2637}, {10'sd501, 13'sd-3514, 13'sd-2655}},
{{7'sd50, 10'sd373, 11'sd-736}, {11'sd-747, 9'sd-181, 10'sd-419}, {13'sd-2931, 12'sd1213, 11'sd515}},
{{12'sd1407, 12'sd1117, 11'sd873}, {12'sd1587, 12'sd-1457, 8'sd-92}, {13'sd-2245, 11'sd-958, 11'sd905}},
{{12'sd-1674, 7'sd-58, 9'sd177}, {12'sd-1281, 9'sd-157, 11'sd-978}, {12'sd1649, 13'sd-2444, 12'sd-1612}},
{{13'sd-2096, 12'sd1998, 11'sd759}, {12'sd1688, 13'sd-2735, 13'sd-2734}, {6'sd30, 12'sd-1206, 13'sd-2387}},
{{12'sd1961, 12'sd-1493, 9'sd-231}, {11'sd868, 11'sd-832, 10'sd-359}, {11'sd-997, 12'sd1031, 12'sd1796}},
{{13'sd-2143, 11'sd-701, 11'sd996}, {9'sd-209, 12'sd-1694, 13'sd-2105}, {13'sd-3355, 12'sd2006, 12'sd1461}},
{{12'sd-1685, 9'sd237, 12'sd1436}, {9'sd-232, 9'sd-158, 13'sd2717}, {13'sd2629, 13'sd2537, 11'sd559}},
{{13'sd2541, 13'sd2440, 10'sd264}, {13'sd-2424, 9'sd-246, 12'sd1745}, {13'sd2061, 12'sd-1364, 12'sd-1844}},
{{11'sd721, 12'sd1125, 12'sd1364}, {12'sd1840, 12'sd-1835, 13'sd-2350}, {12'sd1505, 12'sd1418, 13'sd2547}},
{{11'sd-736, 11'sd-867, 11'sd558}, {8'sd107, 12'sd1310, 11'sd574}, {10'sd343, 11'sd923, 13'sd2063}},
{{12'sd-1321, 13'sd-2160, 13'sd2510}, {12'sd1238, 12'sd1057, 12'sd-1491}, {13'sd-3143, 12'sd-1572, 12'sd1594}},
{{11'sd-534, 12'sd1553, 12'sd1577}, {12'sd-1166, 11'sd834, 13'sd-2336}, {13'sd2063, 12'sd-1276, 12'sd1774}},
{{11'sd-900, 11'sd901, 11'sd-734}, {12'sd-1824, 12'sd1773, 12'sd1683}, {13'sd2382, 13'sd2466, 12'sd1216}},
{{11'sd-857, 13'sd-2077, 8'sd-82}, {9'sd209, 12'sd-1540, 13'sd2495}, {13'sd-2786, 12'sd-1766, 12'sd-1582}},
{{11'sd-976, 11'sd-684, 13'sd-2124}, {13'sd-2054, 11'sd856, 10'sd-407}, {12'sd1578, 11'sd-522, 11'sd567}},
{{12'sd1508, 11'sd916, 12'sd-1389}, {12'sd-1574, 10'sd427, 13'sd-2156}, {13'sd2686, 11'sd792, 8'sd101}},
{{12'sd1894, 11'sd641, 13'sd2163}, {13'sd-3366, 13'sd-3162, 12'sd-1881}, {10'sd-463, 13'sd-2117, 6'sd23}},
{{13'sd2909, 12'sd1165, 11'sd-882}, {13'sd2501, 11'sd674, 12'sd-1165}, {10'sd-321, 12'sd1459, 12'sd1262}},
{{11'sd-659, 13'sd-2694, 12'sd1170}, {7'sd-35, 11'sd866, 10'sd-349}, {13'sd-2448, 12'sd1925, 9'sd169}},
{{12'sd-1076, 11'sd814, 12'sd-1617}, {12'sd1692, 13'sd2242, 13'sd2135}, {13'sd-2543, 12'sd1196, 11'sd-956}},
{{7'sd-46, 12'sd-1289, 12'sd1208}, {13'sd2161, 12'sd1152, 8'sd-91}, {12'sd-1265, 9'sd-132, 12'sd-1657}},
{{12'sd-1520, 13'sd2640, 11'sd1020}, {11'sd-651, 13'sd2752, 11'sd-608}, {11'sd-723, 13'sd-2679, 12'sd1718}},
{{11'sd-1016, 13'sd2467, 12'sd-1144}, {12'sd1207, 12'sd-1863, 11'sd783}, {13'sd2110, 10'sd-292, 10'sd298}},
{{10'sd370, 12'sd-1276, 12'sd1990}, {11'sd791, 11'sd954, 13'sd-2256}, {12'sd1719, 12'sd1508, 12'sd-1109}},
{{8'sd108, 13'sd2438, 8'sd-116}, {5'sd-8, 11'sd-630, 12'sd-1267}, {13'sd2643, 13'sd-2140, 12'sd-1473}},
{{12'sd-1202, 12'sd1214, 12'sd1170}, {11'sd-986, 13'sd-2817, 10'sd309}, {13'sd2724, 11'sd-618, 8'sd-78}},
{{12'sd1407, 9'sd145, 11'sd-670}, {13'sd2788, 13'sd2381, 11'sd-622}, {12'sd-1400, 11'sd-906, 13'sd-2366}},
{{13'sd2262, 11'sd-649, 8'sd98}, {10'sd-272, 11'sd939, 8'sd-82}, {12'sd-1288, 13'sd2203, 8'sd-69}},
{{12'sd-1029, 12'sd1976, 13'sd2055}, {11'sd-535, 12'sd1153, 12'sd1277}, {12'sd-1529, 13'sd3477, 10'sd-341}},
{{13'sd-2064, 12'sd1656, 12'sd1627}, {10'sd451, 13'sd-2495, 10'sd491}, {11'sd1012, 12'sd-1071, 8'sd70}},
{{11'sd787, 12'sd1446, 11'sd616}, {10'sd-352, 13'sd-2807, 12'sd1678}, {10'sd-359, 13'sd2431, 6'sd31}},
{{10'sd-420, 11'sd-828, 12'sd-1065}, {11'sd899, 13'sd2556, 12'sd1668}, {11'sd-918, 12'sd-1356, 12'sd1311}},
{{12'sd1957, 11'sd-1016, 10'sd501}, {11'sd-864, 11'sd-524, 11'sd741}, {13'sd2258, 8'sd116, 11'sd756}},
{{13'sd2134, 11'sd-725, 12'sd-1711}, {12'sd2030, 12'sd-1941, 10'sd495}, {10'sd-261, 12'sd1777, 10'sd-438}},
{{10'sd-419, 8'sd-85, 12'sd1171}, {10'sd-510, 12'sd1742, 12'sd-1475}, {8'sd-75, 12'sd-1617, 9'sd-252}},
{{11'sd-693, 12'sd-1086, 7'sd-43}, {11'sd888, 8'sd-94, 9'sd138}, {12'sd-1654, 11'sd-874, 11'sd953}},
{{10'sd349, 12'sd1806, 12'sd-1461}, {13'sd2118, 12'sd-1199, 13'sd-2357}, {12'sd-1747, 13'sd2407, 11'sd684}},
{{12'sd1321, 12'sd-1684, 13'sd-2204}, {9'sd-151, 11'sd-513, 13'sd-2835}, {10'sd-332, 13'sd2084, 12'sd1026}},
{{12'sd-1101, 13'sd-2628, 12'sd-1733}, {10'sd-381, 13'sd3209, 13'sd2608}, {13'sd3017, 12'sd-1650, 8'sd-126}},
{{10'sd477, 13'sd-2403, 13'sd-2323}, {12'sd1637, 13'sd2247, 12'sd-1312}, {11'sd-737, 12'sd-1606, 12'sd1339}},
{{12'sd-1818, 10'sd-467, 12'sd-1198}, {12'sd-1112, 13'sd2088, 12'sd1165}, {12'sd-1418, 11'sd611, 11'sd817}},
{{8'sd-91, 12'sd1694, 12'sd-1199}, {12'sd1933, 12'sd-1479, 11'sd-600}, {12'sd-1967, 8'sd-126, 10'sd-483}},
{{13'sd2505, 10'sd-269, 13'sd2332}, {13'sd-2954, 13'sd-2401, 13'sd2524}, {12'sd-1780, 7'sd-38, 13'sd-2480}},
{{9'sd162, 12'sd-1538, 11'sd-901}, {12'sd-1049, 12'sd1647, 13'sd2311}, {13'sd2555, 12'sd1923, 13'sd2311}},
{{12'sd-1955, 11'sd-753, 10'sd368}, {7'sd55, 13'sd3003, 13'sd-2632}, {13'sd4085, 11'sd-836, 10'sd-308}},
{{13'sd2349, 13'sd-2069, 13'sd-2109}, {10'sd311, 13'sd2528, 12'sd-1787}, {11'sd-595, 11'sd780, 8'sd-122}},
{{10'sd292, 13'sd-2442, 11'sd-796}, {13'sd-2592, 12'sd-1093, 11'sd561}, {12'sd1861, 12'sd-1318, 12'sd-1288}},
{{7'sd56, 13'sd-2741, 12'sd-1333}, {12'sd2020, 10'sd-260, 6'sd-21}, {13'sd2161, 11'sd778, 13'sd2975}},
{{7'sd56, 13'sd-2093, 13'sd-2202}, {8'sd-75, 13'sd-2808, 13'sd2451}, {11'sd598, 11'sd579, 11'sd-962}},
{{13'sd2651, 11'sd-631, 12'sd1123}, {9'sd-199, 11'sd539, 13'sd2130}, {12'sd-1542, 13'sd-2494, 10'sd-470}},
{{12'sd-1413, 11'sd615, 11'sd-1003}, {9'sd251, 13'sd2821, 12'sd1382}, {13'sd3329, 12'sd-1671, 10'sd505}},
{{11'sd-774, 12'sd1107, 13'sd-2323}, {11'sd1007, 12'sd-1589, 12'sd-1157}, {13'sd-2896, 10'sd-461, 13'sd-2569}},
{{11'sd618, 13'sd3058, 11'sd799}, {13'sd2361, 11'sd-645, 7'sd53}, {12'sd1998, 13'sd-2813, 6'sd-16}},
{{13'sd-2270, 11'sd547, 13'sd2747}, {11'sd895, 13'sd-2349, 10'sd-275}, {13'sd-2272, 12'sd1161, 12'sd-1222}},
{{12'sd2033, 12'sd-1036, 13'sd2587}, {12'sd1497, 13'sd-2680, 10'sd-493}, {13'sd-3018, 11'sd891, 11'sd804}},
{{13'sd-2311, 11'sd-1007, 13'sd-2470}, {13'sd-2641, 12'sd1600, 11'sd-974}, {11'sd-683, 12'sd1064, 10'sd302}}},
{
{{14'sd4331, 13'sd3913, 12'sd1574}, {13'sd2913, 13'sd3123, 13'sd3255}, {13'sd-2689, 14'sd-4236, 12'sd1156}},
{{10'sd506, 13'sd2149, 13'sd-2395}, {12'sd1068, 12'sd-1977, 12'sd-1148}, {12'sd-1856, 11'sd556, 12'sd-1683}},
{{12'sd1181, 13'sd3433, 12'sd1618}, {13'sd2230, 12'sd1601, 12'sd-1314}, {13'sd-3108, 10'sd437, 13'sd-2314}},
{{12'sd-1496, 13'sd-2119, 12'sd-1813}, {13'sd-2317, 12'sd-1353, 13'sd2308}, {8'sd-126, 12'sd1434, 12'sd-1529}},
{{13'sd2277, 11'sd704, 13'sd2222}, {13'sd3088, 10'sd-462, 11'sd-909}, {13'sd2997, 13'sd-3030, 11'sd-923}},
{{10'sd-309, 12'sd-1202, 11'sd-833}, {12'sd1396, 8'sd70, 13'sd2050}, {11'sd-963, 12'sd-1190, 14'sd4144}},
{{10'sd-324, 12'sd1101, 12'sd1189}, {11'sd662, 10'sd-490, 12'sd-1896}, {13'sd2662, 12'sd1439, 12'sd1883}},
{{11'sd-791, 13'sd-2436, 11'sd-558}, {12'sd1835, 13'sd2549, 9'sd-143}, {12'sd1496, 13'sd2423, 11'sd993}},
{{9'sd-213, 12'sd-1088, 13'sd-2469}, {12'sd-2011, 11'sd-914, 12'sd1315}, {11'sd-736, 8'sd106, 10'sd-283}},
{{4'sd6, 12'sd1369, 12'sd1971}, {13'sd3227, 12'sd1987, 8'sd87}, {13'sd-2256, 13'sd3897, 12'sd1796}},
{{13'sd3562, 11'sd-724, 11'sd895}, {10'sd-484, 13'sd-2616, 13'sd2449}, {13'sd4074, 13'sd2998, 13'sd3547}},
{{12'sd1274, 11'sd-992, 11'sd-932}, {13'sd3297, 11'sd655, 12'sd1523}, {13'sd-2388, 11'sd-991, 12'sd-1695}},
{{14'sd-4564, 13'sd-3554, 14'sd-4208}, {12'sd-1544, 13'sd-2125, 12'sd-1648}, {13'sd3447, 12'sd1181, 13'sd2956}},
{{11'sd-861, 9'sd187, 13'sd-2117}, {11'sd798, 13'sd-2433, 13'sd2374}, {12'sd1742, 12'sd-1902, 13'sd3104}},
{{10'sd-350, 12'sd-1560, 13'sd-2205}, {11'sd727, 13'sd-2924, 13'sd-2627}, {11'sd-873, 11'sd-608, 12'sd-1560}},
{{9'sd238, 10'sd-443, 11'sd530}, {11'sd903, 12'sd-1953, 12'sd1987}, {13'sd3268, 13'sd3318, 13'sd3263}},
{{12'sd1863, 10'sd385, 13'sd-3013}, {11'sd-979, 12'sd1446, 11'sd-616}, {11'sd553, 14'sd4470, 7'sd48}},
{{13'sd2992, 10'sd310, 10'sd256}, {12'sd-1249, 10'sd485, 13'sd-2543}, {13'sd-2108, 8'sd-96, 6'sd30}},
{{11'sd883, 11'sd-581, 11'sd659}, {12'sd-1880, 11'sd549, 13'sd2491}, {13'sd-2422, 12'sd-1201, 12'sd1161}},
{{13'sd2260, 13'sd-2761, 11'sd-586}, {13'sd2586, 9'sd-239, 10'sd481}, {13'sd3421, 13'sd4047, 9'sd164}},
{{12'sd-1393, 13'sd2175, 10'sd377}, {13'sd2782, 11'sd-523, 10'sd-506}, {9'sd-253, 7'sd-63, 12'sd1938}},
{{13'sd-3526, 12'sd1522, 12'sd-1285}, {11'sd722, 12'sd-1346, 11'sd-847}, {13'sd3390, 12'sd1117, 12'sd-1415}},
{{11'sd651, 12'sd1540, 11'sd802}, {13'sd2836, 12'sd1100, 13'sd-2390}, {13'sd-2150, 10'sd299, 5'sd12}},
{{13'sd-2584, 13'sd-2477, 11'sd-862}, {12'sd-1056, 13'sd-2124, 13'sd2501}, {11'sd-759, 9'sd206, 12'sd-1194}},
{{11'sd933, 9'sd130, 11'sd-638}, {13'sd2368, 13'sd3118, 12'sd1283}, {13'sd-2288, 14'sd-4418, 13'sd-2573}},
{{12'sd-1786, 11'sd-618, 13'sd-2060}, {12'sd1148, 13'sd-2557, 12'sd1540}, {13'sd-2215, 11'sd-967, 10'sd428}},
{{9'sd-239, 13'sd-3037, 12'sd1582}, {10'sd-431, 12'sd1907, 13'sd2213}, {12'sd1704, 13'sd2061, 10'sd-294}},
{{12'sd-1715, 9'sd-156, 10'sd463}, {10'sd-450, 7'sd-32, 11'sd-689}, {12'sd-1137, 11'sd-851, 11'sd-675}},
{{12'sd-1856, 11'sd-665, 11'sd652}, {11'sd514, 8'sd114, 8'sd-93}, {13'sd2864, 12'sd1409, 7'sd-59}},
{{10'sd-265, 12'sd1782, 11'sd-874}, {12'sd1849, 12'sd-1421, 12'sd-1658}, {13'sd3426, 12'sd-1806, 10'sd-262}},
{{12'sd-1747, 12'sd1818, 12'sd-1463}, {13'sd-2205, 13'sd2169, 12'sd-1143}, {11'sd757, 13'sd3429, 12'sd-1300}},
{{11'sd978, 11'sd991, 9'sd133}, {12'sd1595, 12'sd2014, 11'sd953}, {13'sd2113, 12'sd1658, 9'sd177}},
{{13'sd2202, 13'sd2972, 12'sd1860}, {13'sd2659, 13'sd3759, 13'sd-2181}, {12'sd1746, 12'sd1692, 13'sd-3157}},
{{13'sd-2254, 12'sd1806, 11'sd642}, {13'sd-2833, 12'sd-1459, 11'sd-741}, {12'sd1380, 13'sd2110, 11'sd626}},
{{14'sd4118, 12'sd-1066, 11'sd1015}, {13'sd2937, 12'sd2043, 13'sd2967}, {13'sd-2052, 13'sd-3055, 12'sd1526}},
{{13'sd2586, 12'sd-1297, 10'sd-354}, {10'sd-481, 10'sd-349, 13'sd3000}, {12'sd-1913, 9'sd-224, 13'sd2584}},
{{12'sd1024, 13'sd-2329, 9'sd153}, {10'sd-494, 12'sd1866, 13'sd-3050}, {9'sd250, 13'sd-2368, 11'sd-664}},
{{8'sd108, 13'sd-2431, 12'sd1957}, {13'sd3133, 13'sd2469, 10'sd-282}, {12'sd-1648, 13'sd-2528, 13'sd-3480}},
{{13'sd2653, 10'sd-306, 4'sd-5}, {9'sd142, 12'sd-1128, 13'sd-2486}, {14'sd4599, 13'sd2682, 13'sd-2146}},
{{11'sd-540, 13'sd-2751, 4'sd5}, {12'sd1321, 9'sd-214, 11'sd542}, {12'sd-1960, 12'sd-1100, 11'sd-857}},
{{12'sd1212, 10'sd-482, 12'sd1299}, {11'sd821, 13'sd2474, 13'sd-3357}, {10'sd-322, 12'sd1057, 12'sd1845}},
{{13'sd-2847, 13'sd2427, 12'sd1963}, {12'sd-2021, 11'sd-532, 13'sd2371}, {13'sd-3334, 8'sd92, 13'sd-3430}},
{{12'sd1871, 13'sd-2925, 13'sd-2153}, {13'sd2416, 9'sd-136, 9'sd190}, {13'sd2806, 12'sd1111, 12'sd1027}},
{{11'sd-1005, 10'sd-434, 11'sd-749}, {12'sd-1055, 12'sd-1997, 12'sd1291}, {13'sd-2332, 12'sd1583, 13'sd2491}},
{{13'sd-2357, 12'sd-1397, 9'sd-237}, {12'sd1187, 13'sd-2915, 13'sd-2310}, {13'sd2740, 13'sd2171, 13'sd-2464}},
{{13'sd-2607, 12'sd1336, 10'sd346}, {11'sd-721, 13'sd-2465, 13'sd-2495}, {11'sd524, 13'sd-2569, 14'sd-4327}},
{{12'sd1927, 13'sd3129, 11'sd-713}, {12'sd-1281, 11'sd-905, 13'sd-2842}, {12'sd-1308, 9'sd247, 12'sd-1381}},
{{11'sd575, 12'sd1715, 12'sd1956}, {12'sd-1400, 12'sd-1452, 13'sd2351}, {13'sd-2353, 12'sd1179, 12'sd-1940}},
{{11'sd-531, 12'sd1350, 10'sd445}, {11'sd-647, 10'sd-450, 13'sd2938}, {12'sd-1992, 13'sd-3193, 12'sd1250}},
{{12'sd-1071, 13'sd-2644, 13'sd-2537}, {12'sd-1283, 13'sd2410, 11'sd-629}, {13'sd2187, 10'sd500, 12'sd-1255}},
{{11'sd572, 13'sd-2865, 11'sd-516}, {12'sd1582, 11'sd951, 13'sd-2429}, {12'sd1737, 12'sd1363, 12'sd-1858}},
{{12'sd-1110, 11'sd-821, 12'sd1465}, {11'sd-556, 11'sd694, 12'sd-1354}, {11'sd705, 13'sd-2197, 13'sd2365}},
{{13'sd-2529, 13'sd2321, 11'sd-888}, {12'sd-1047, 12'sd1476, 13'sd-2782}, {12'sd1127, 13'sd-3163, 13'sd-3280}},
{{11'sd582, 11'sd1003, 12'sd1267}, {12'sd1342, 6'sd-27, 11'sd850}, {13'sd2607, 12'sd-1133, 11'sd827}},
{{11'sd826, 12'sd1935, 10'sd-393}, {10'sd-347, 13'sd2367, 11'sd932}, {9'sd-154, 11'sd562, 12'sd1131}},
{{12'sd-1584, 13'sd-2768, 12'sd-1744}, {13'sd-2266, 13'sd-2098, 12'sd1418}, {13'sd-2079, 13'sd2100, 13'sd-2136}},
{{12'sd-1735, 13'sd-3332, 13'sd-2077}, {12'sd-1622, 12'sd1157, 12'sd1076}, {10'sd-390, 12'sd-1809, 11'sd634}},
{{12'sd-1528, 12'sd-1638, 11'sd782}, {14'sd-4567, 12'sd1511, 13'sd-2477}, {14'sd-7109, 12'sd1517, 13'sd2714}},
{{13'sd3576, 6'sd-31, 10'sd357}, {11'sd803, 13'sd-2453, 12'sd1039}, {13'sd2139, 13'sd3275, 14'sd5764}},
{{13'sd-2935, 11'sd-1022, 11'sd786}, {12'sd1343, 9'sd-131, 12'sd-1968}, {11'sd943, 11'sd965, 12'sd-1790}},
{{13'sd2559, 13'sd2232, 11'sd593}, {13'sd2108, 11'sd640, 11'sd688}, {12'sd1765, 12'sd1664, 10'sd307}},
{{12'sd-1793, 10'sd-405, 13'sd2127}, {11'sd-858, 11'sd-569, 11'sd-992}, {12'sd-1189, 12'sd1990, 12'sd1516}},
{{13'sd-2102, 7'sd52, 13'sd-2759}, {12'sd-1309, 11'sd-804, 13'sd-2870}, {10'sd-325, 12'sd1533, 10'sd306}},
{{11'sd-850, 9'sd216, 12'sd-1298}, {11'sd908, 13'sd2606, 10'sd-312}, {12'sd1378, 13'sd-3917, 12'sd1581}}},
{
{{13'sd2072, 11'sd738, 12'sd-1260}, {11'sd853, 10'sd-425, 12'sd1243}, {13'sd2250, 13'sd2186, 13'sd2129}},
{{12'sd1727, 13'sd-2193, 13'sd-2943}, {12'sd1788, 12'sd1650, 11'sd-637}, {12'sd-1682, 13'sd3006, 12'sd1572}},
{{14'sd4106, 13'sd3691, 9'sd205}, {10'sd-349, 8'sd80, 13'sd2065}, {11'sd-564, 8'sd-82, 13'sd-2315}},
{{13'sd-2741, 11'sd-785, 11'sd767}, {12'sd2009, 12'sd-1350, 12'sd-1536}, {11'sd1020, 12'sd1063, 13'sd-2416}},
{{12'sd1718, 12'sd-1919, 12'sd1820}, {11'sd-750, 13'sd-3255, 12'sd1394}, {12'sd-1737, 7'sd-44, 12'sd1184}},
{{12'sd1924, 11'sd681, 7'sd-39}, {12'sd1528, 12'sd1380, 9'sd239}, {13'sd2333, 9'sd208, 9'sd254}},
{{12'sd1465, 12'sd-1475, 11'sd-854}, {10'sd-357, 11'sd-815, 12'sd1556}, {12'sd-1773, 12'sd-1123, 11'sd684}},
{{13'sd-2075, 8'sd65, 12'sd1055}, {12'sd-1642, 12'sd1211, 12'sd-1724}, {13'sd3405, 11'sd-750, 12'sd1978}},
{{7'sd-53, 11'sd-937, 12'sd1397}, {9'sd232, 13'sd2322, 8'sd-73}, {10'sd-358, 13'sd3059, 11'sd574}},
{{10'sd-489, 10'sd410, 13'sd-3093}, {13'sd2455, 10'sd-323, 12'sd1282}, {12'sd-1101, 7'sd47, 12'sd1191}},
{{13'sd-3744, 13'sd-3085, 11'sd-604}, {12'sd-1030, 11'sd1000, 11'sd-613}, {13'sd-2339, 13'sd-2769, 13'sd2069}},
{{13'sd-2446, 13'sd-2472, 10'sd-421}, {12'sd-1074, 13'sd-2345, 13'sd-2441}, {11'sd-527, 11'sd742, 12'sd1085}},
{{7'sd-62, 12'sd-1550, 12'sd-1205}, {11'sd-544, 10'sd290, 13'sd-2904}, {12'sd1623, 13'sd2554, 13'sd-2894}},
{{12'sd1947, 12'sd-1276, 11'sd-640}, {11'sd-693, 12'sd-1160, 12'sd-2004}, {13'sd2599, 10'sd-367, 12'sd-2043}},
{{12'sd1515, 10'sd-320, 13'sd-2090}, {11'sd554, 12'sd1192, 12'sd-1576}, {13'sd2098, 11'sd725, 11'sd904}},
{{11'sd-749, 13'sd-2873, 13'sd-2824}, {12'sd-1216, 11'sd825, 12'sd1045}, {13'sd3082, 12'sd-1701, 11'sd-933}},
{{7'sd37, 13'sd-2665, 12'sd1088}, {12'sd-1660, 12'sd-1109, 12'sd1128}, {11'sd986, 12'sd-1065, 13'sd-2525}},
{{13'sd2610, 14'sd4172, 8'sd-118}, {12'sd1989, 12'sd1802, 12'sd1103}, {13'sd-2509, 12'sd-1287, 13'sd-3095}},
{{12'sd1413, 12'sd-1611, 10'sd364}, {12'sd-1186, 13'sd-2807, 11'sd994}, {11'sd761, 12'sd-1995, 12'sd-1291}},
{{12'sd1078, 12'sd-1550, 11'sd-597}, {10'sd-495, 13'sd-2051, 13'sd-2845}, {12'sd-1523, 13'sd-2602, 12'sd-1984}},
{{9'sd150, 11'sd864, 10'sd-485}, {10'sd412, 8'sd-100, 11'sd-694}, {13'sd-2549, 12'sd-1278, 12'sd-1800}},
{{12'sd-1269, 11'sd-825, 13'sd-2311}, {10'sd274, 13'sd-3488, 10'sd302}, {11'sd-788, 11'sd1018, 13'sd2400}},
{{12'sd1068, 10'sd-362, 11'sd-984}, {11'sd698, 13'sd3052, 12'sd1735}, {10'sd285, 13'sd-2496, 12'sd1949}},
{{12'sd-1620, 12'sd-2040, 13'sd2946}, {12'sd-1557, 8'sd71, 13'sd2054}, {13'sd-2485, 10'sd-389, 11'sd979}},
{{13'sd4061, 12'sd1703, 11'sd-840}, {13'sd3748, 13'sd3517, 11'sd881}, {13'sd3380, 11'sd-832, 9'sd134}},
{{12'sd1737, 13'sd-2713, 13'sd2309}, {13'sd-2060, 13'sd-2723, 13'sd2388}, {10'sd399, 12'sd1059, 12'sd-1449}},
{{13'sd2442, 11'sd-682, 13'sd2263}, {9'sd157, 7'sd44, 12'sd-1441}, {10'sd281, 10'sd-351, 9'sd-148}},
{{10'sd354, 9'sd-168, 12'sd1844}, {11'sd-536, 12'sd1140, 11'sd-668}, {12'sd-1976, 12'sd-1611, 11'sd1008}},
{{9'sd-234, 12'sd-1043, 12'sd1496}, {13'sd-2777, 7'sd59, 8'sd125}, {12'sd2023, 9'sd210, 13'sd2188}},
{{11'sd699, 11'sd-939, 11'sd-852}, {10'sd497, 12'sd-1969, 13'sd2094}, {11'sd555, 12'sd1617, 12'sd1684}},
{{13'sd-2284, 13'sd-2268, 12'sd-1811}, {7'sd33, 13'sd-2349, 12'sd-1297}, {10'sd-413, 11'sd-571, 12'sd-1620}},
{{13'sd-2568, 12'sd1812, 12'sd-1432}, {9'sd214, 12'sd-1569, 12'sd-1187}, {11'sd527, 12'sd-1762, 10'sd-486}},
{{12'sd-1192, 13'sd2139, 13'sd2073}, {13'sd2095, 13'sd-2254, 10'sd348}, {11'sd581, 13'sd-2850, 9'sd187}},
{{12'sd-1041, 12'sd-2031, 7'sd-33}, {12'sd-1068, 12'sd1490, 10'sd-406}, {13'sd2430, 10'sd-456, 12'sd-1108}},
{{13'sd-3335, 13'sd2283, 12'sd-1552}, {9'sd-170, 13'sd2251, 12'sd2012}, {11'sd968, 12'sd1179, 12'sd1733}},
{{11'sd985, 12'sd1988, 13'sd2337}, {11'sd-807, 13'sd2386, 13'sd2143}, {13'sd2310, 11'sd581, 12'sd1757}},
{{12'sd1750, 13'sd3484, 13'sd2528}, {13'sd2186, 12'sd-1712, 12'sd1150}, {10'sd-329, 12'sd1326, 8'sd103}},
{{12'sd1305, 13'sd-3015, 7'sd62}, {10'sd-419, 11'sd-975, 12'sd1751}, {13'sd2282, 12'sd-1911, 12'sd1050}},
{{12'sd-1326, 7'sd-61, 13'sd-3150}, {11'sd692, 12'sd-1946, 13'sd-3223}, {12'sd-1179, 11'sd1003, 11'sd841}},
{{12'sd1501, 12'sd-1262, 11'sd994}, {10'sd-334, 12'sd-1447, 11'sd711}, {10'sd275, 8'sd-73, 9'sd220}},
{{10'sd291, 12'sd1816, 12'sd-1923}, {11'sd847, 9'sd204, 12'sd1525}, {11'sd-622, 11'sd974, 12'sd-1777}},
{{11'sd-954, 13'sd-2617, 12'sd1087}, {13'sd2505, 13'sd2348, 12'sd1417}, {13'sd-2117, 9'sd-129, 12'sd1805}},
{{12'sd1414, 13'sd-2232, 8'sd-124}, {12'sd-1773, 7'sd42, 12'sd-1640}, {11'sd-617, 12'sd1929, 10'sd464}},
{{12'sd1138, 12'sd1621, 12'sd-1960}, {12'sd-1772, 13'sd-2679, 11'sd-685}, {11'sd-784, 8'sd-96, 11'sd-958}},
{{11'sd-566, 11'sd695, 12'sd1390}, {13'sd2195, 13'sd2190, 12'sd-1751}, {12'sd1305, 12'sd1944, 12'sd-1778}},
{{11'sd998, 13'sd-2088, 12'sd-1526}, {12'sd-1645, 11'sd-964, 8'sd-93}, {13'sd2345, 11'sd975, 11'sd647}},
{{13'sd2171, 13'sd-2119, 11'sd-805}, {10'sd-471, 12'sd-1884, 11'sd-646}, {11'sd-735, 11'sd-902, 7'sd-49}},
{{12'sd1444, 12'sd-1295, 12'sd-1487}, {10'sd-326, 12'sd-1752, 12'sd1187}, {11'sd1016, 13'sd-2100, 13'sd2619}},
{{12'sd1402, 13'sd-2420, 12'sd-1816}, {11'sd838, 10'sd-272, 12'sd-1267}, {10'sd-293, 10'sd-410, 13'sd2814}},
{{10'sd354, 13'sd-2155, 13'sd2674}, {11'sd-582, 11'sd831, 13'sd2487}, {12'sd1391, 11'sd-525, 13'sd2352}},
{{12'sd-1931, 8'sd76, 9'sd-151}, {10'sd368, 12'sd-1204, 12'sd1617}, {11'sd927, 11'sd-543, 11'sd-745}},
{{10'sd359, 10'sd304, 12'sd2015}, {12'sd1140, 12'sd1992, 13'sd-2090}, {13'sd-2544, 12'sd-1772, 13'sd-2442}},
{{12'sd1932, 10'sd-261, 11'sd-743}, {12'sd-1565, 9'sd-147, 13'sd3432}, {12'sd1415, 11'sd572, 11'sd705}},
{{11'sd-974, 11'sd871, 10'sd-410}, {12'sd1364, 12'sd-1515, 10'sd-498}, {13'sd2097, 12'sd1398, 11'sd-689}},
{{12'sd1727, 13'sd2654, 11'sd-724}, {12'sd-1063, 12'sd1157, 12'sd1471}, {12'sd1141, 12'sd-1567, 12'sd1868}},
{{10'sd408, 12'sd-1762, 13'sd2805}, {11'sd-723, 13'sd3006, 9'sd-134}, {12'sd1381, 11'sd-748, 12'sd-2031}},
{{10'sd-511, 12'sd-1130, 12'sd-1903}, {11'sd-531, 11'sd626, 11'sd789}, {13'sd-2697, 12'sd1733, 13'sd2597}},
{{13'sd-2759, 10'sd-449, 12'sd-1324}, {12'sd1676, 11'sd565, 13'sd2149}, {12'sd1239, 9'sd150, 13'sd-2305}},
{{13'sd2510, 12'sd1837, 12'sd1434}, {13'sd-2455, 7'sd42, 11'sd770}, {12'sd-1452, 12'sd-1232, 12'sd-1375}},
{{13'sd-2691, 13'sd-2762, 12'sd-1729}, {12'sd1768, 12'sd1542, 10'sd462}, {12'sd1362, 13'sd-2122, 13'sd-2432}},
{{11'sd695, 7'sd-63, 13'sd2610}, {11'sd743, 12'sd1817, 12'sd-1429}, {13'sd2794, 13'sd2401, 11'sd-938}},
{{12'sd-1231, 13'sd-2853, 12'sd1291}, {12'sd1620, 13'sd-2269, 11'sd602}, {13'sd2525, 11'sd893, 8'sd-115}},
{{9'sd144, 11'sd587, 11'sd-1016}, {12'sd-1378, 12'sd1116, 9'sd-232}, {11'sd-903, 12'sd-1185, 10'sd-310}},
{{12'sd-1685, 13'sd2450, 11'sd-810}, {8'sd-68, 11'sd-851, 12'sd-1523}, {11'sd-578, 13'sd2089, 12'sd-1897}}},
{
{{12'sd1283, 12'sd-1441, 6'sd27}, {11'sd707, 12'sd-1682, 13'sd-2322}, {13'sd-2735, 13'sd-2828, 13'sd-2287}},
{{13'sd-2768, 12'sd-1905, 12'sd-1665}, {12'sd1403, 10'sd-373, 11'sd-1002}, {9'sd-148, 12'sd1480, 11'sd1023}},
{{12'sd1979, 13'sd-3605, 11'sd-741}, {10'sd-290, 11'sd980, 11'sd959}, {13'sd3784, 12'sd1949, 12'sd-1655}},
{{8'sd-99, 11'sd706, 11'sd-597}, {12'sd-1672, 12'sd1465, 12'sd-1290}, {12'sd-1539, 12'sd1047, 12'sd-1369}},
{{13'sd2705, 11'sd-626, 12'sd1606}, {13'sd3286, 10'sd360, 12'sd-1682}, {13'sd-2921, 12'sd-1152, 13'sd-2226}},
{{13'sd-2805, 10'sd-416, 12'sd1024}, {11'sd-821, 10'sd484, 13'sd2096}, {11'sd916, 12'sd1491, 8'sd106}},
{{14'sd4618, 13'sd2598, 14'sd5124}, {12'sd-1162, 11'sd-540, 12'sd1911}, {13'sd-2385, 13'sd2173, 10'sd290}},
{{14'sd4203, 11'sd775, 11'sd-971}, {12'sd1696, 11'sd-929, 13'sd-2855}, {13'sd3651, 12'sd-1838, 13'sd-3922}},
{{12'sd-1211, 13'sd-3030, 13'sd-4069}, {13'sd2166, 12'sd1613, 12'sd-1527}, {13'sd3689, 11'sd-979, 12'sd1760}},
{{10'sd474, 12'sd-1035, 10'sd333}, {11'sd-524, 13'sd2055, 12'sd-1118}, {11'sd-1017, 12'sd1392, 13'sd-3217}},
{{13'sd-2541, 5'sd9, 14'sd5075}, {12'sd1357, 13'sd3181, 13'sd3815}, {13'sd3786, 14'sd5260, 14'sd5118}},
{{13'sd2160, 12'sd1494, 13'sd2922}, {12'sd-1484, 12'sd1144, 9'sd143}, {11'sd-578, 12'sd1889, 10'sd-331}},
{{12'sd-1539, 10'sd369, 13'sd-2057}, {11'sd849, 5'sd14, 13'sd-3509}, {12'sd1663, 11'sd-666, 12'sd-1186}},
{{11'sd548, 11'sd726, 12'sd-1655}, {12'sd-1731, 11'sd660, 13'sd-2795}, {12'sd-1079, 11'sd-732, 13'sd2197}},
{{11'sd780, 12'sd1430, 8'sd-121}, {12'sd1188, 12'sd-1261, 12'sd-1586}, {13'sd-2765, 11'sd-937, 10'sd-314}},
{{13'sd2729, 12'sd1308, 13'sd-2400}, {13'sd2666, 10'sd-295, 11'sd859}, {13'sd2457, 12'sd1158, 12'sd1446}},
{{13'sd2121, 12'sd-1285, 13'sd2823}, {12'sd1714, 10'sd301, 10'sd-338}, {11'sd560, 13'sd-2535, 12'sd1901}},
{{13'sd2873, 13'sd-2533, 12'sd-1699}, {12'sd1105, 13'sd2211, 13'sd-2439}, {9'sd230, 11'sd570, 14'sd-4580}},
{{14'sd4100, 9'sd179, 12'sd-1504}, {11'sd-761, 12'sd-1105, 13'sd-2505}, {12'sd1817, 12'sd-1896, 13'sd-2243}},
{{12'sd1656, 12'sd-1513, 14'sd-4104}, {9'sd218, 11'sd618, 13'sd-2387}, {13'sd-2209, 11'sd-753, 12'sd1527}},
{{13'sd-3998, 14'sd-4115, 14'sd-4109}, {11'sd-623, 11'sd-817, 12'sd-2013}, {13'sd2137, 8'sd-69, 12'sd-1516}},
{{13'sd-3899, 12'sd1425, 14'sd5408}, {14'sd-4817, 13'sd-2821, 10'sd382}, {13'sd-3948, 11'sd-589, 12'sd1931}},
{{10'sd366, 11'sd-629, 12'sd-1345}, {13'sd-2254, 9'sd-202, 13'sd-2563}, {13'sd-2066, 12'sd1115, 11'sd-919}},
{{12'sd-1354, 10'sd478, 12'sd-1674}, {11'sd698, 12'sd-1299, 13'sd-2451}, {13'sd2400, 10'sd446, 13'sd-2165}},
{{13'sd-2352, 10'sd-410, 6'sd18}, {12'sd1476, 8'sd-106, 13'sd-2574}, {12'sd1254, 11'sd521, 13'sd-2532}},
{{12'sd-1114, 12'sd1415, 10'sd-483}, {10'sd-454, 12'sd-1256, 11'sd-798}, {12'sd1807, 12'sd1237, 12'sd1720}},
{{13'sd2995, 13'sd2868, 10'sd401}, {13'sd-2058, 13'sd-2176, 11'sd-997}, {12'sd1960, 12'sd-1510, 12'sd-1034}},
{{7'sd-57, 10'sd296, 11'sd-559}, {13'sd2923, 12'sd-1404, 12'sd-1285}, {11'sd-889, 11'sd-562, 12'sd-1335}},
{{11'sd-589, 11'sd-963, 13'sd3710}, {12'sd-1161, 11'sd-942, 10'sd345}, {13'sd-3762, 13'sd2947, 12'sd1786}},
{{11'sd-778, 11'sd606, 10'sd-260}, {12'sd-1388, 12'sd1504, 13'sd3369}, {13'sd-3211, 13'sd-2473, 11'sd830}},
{{12'sd1681, 12'sd-1623, 6'sd-22}, {11'sd-990, 12'sd1945, 12'sd-1066}, {13'sd-2493, 13'sd2555, 12'sd-1132}},
{{11'sd882, 13'sd2201, 9'sd-213}, {13'sd3218, 13'sd-2086, 11'sd994}, {12'sd1554, 11'sd-836, 12'sd-1353}},
{{11'sd887, 11'sd592, 12'sd1526}, {13'sd2773, 12'sd1743, 10'sd-257}, {11'sd-971, 7'sd-52, 13'sd2634}},
{{11'sd-811, 12'sd1407, 13'sd2356}, {13'sd-3017, 12'sd1076, 12'sd-1178}, {10'sd-418, 12'sd1418, 13'sd2860}},
{{12'sd1708, 12'sd1526, 12'sd-1210}, {12'sd1742, 13'sd2082, 11'sd-556}, {9'sd142, 12'sd-1266, 12'sd-1149}},
{{12'sd-1889, 12'sd-1871, 13'sd2715}, {12'sd-1817, 13'sd-2910, 12'sd1553}, {13'sd2338, 11'sd860, 12'sd1398}},
{{13'sd-3157, 13'sd-2260, 12'sd-1038}, {12'sd-1645, 13'sd2218, 11'sd636}, {10'sd-470, 13'sd2696, 12'sd1489}},
{{11'sd-720, 8'sd127, 10'sd484}, {12'sd1699, 11'sd512, 11'sd915}, {13'sd-2550, 13'sd-3026, 9'sd-239}},
{{13'sd3112, 11'sd-581, 11'sd-566}, {12'sd1257, 10'sd465, 7'sd42}, {12'sd-1454, 13'sd-2892, 13'sd-2927}},
{{14'sd4131, 13'sd2287, 12'sd1336}, {13'sd3149, 7'sd-63, 10'sd-430}, {12'sd1225, 9'sd244, 11'sd922}},
{{11'sd841, 13'sd-3340, 9'sd-165}, {12'sd-1240, 13'sd2479, 12'sd1032}, {12'sd-2024, 11'sd884, 11'sd593}},
{{12'sd1457, 9'sd213, 13'sd2631}, {11'sd-627, 12'sd1748, 10'sd276}, {12'sd1377, 12'sd1322, 13'sd-2322}},
{{11'sd771, 11'sd569, 9'sd-180}, {13'sd2344, 11'sd607, 13'sd-3026}, {12'sd-1923, 11'sd-695, 12'sd-1105}},
{{12'sd1378, 12'sd1423, 12'sd1940}, {10'sd-490, 9'sd231, 11'sd-599}, {12'sd1441, 11'sd-883, 10'sd-260}},
{{12'sd-1101, 4'sd4, 13'sd-3131}, {13'sd-2491, 12'sd1069, 10'sd436}, {9'sd-246, 12'sd1075, 12'sd1617}},
{{13'sd-3306, 13'sd-2080, 12'sd-1174}, {13'sd-2447, 12'sd1268, 10'sd402}, {13'sd2284, 10'sd368, 10'sd341}},
{{11'sd512, 14'sd4272, 13'sd3882}, {9'sd230, 12'sd-1380, 10'sd-400}, {9'sd205, 12'sd-1429, 13'sd-2068}},
{{13'sd-2749, 9'sd-252, 12'sd1689}, {12'sd-1635, 10'sd-464, 12'sd-1615}, {11'sd-878, 9'sd-244, 13'sd2179}},
{{12'sd1989, 10'sd323, 13'sd3119}, {11'sd792, 12'sd-1564, 11'sd-950}, {12'sd-1584, 12'sd1734, 11'sd826}},
{{12'sd1087, 11'sd-710, 12'sd1366}, {12'sd1676, 11'sd-562, 9'sd-226}, {11'sd-732, 12'sd1895, 12'sd-2036}},
{{13'sd2314, 12'sd-1417, 12'sd-1363}, {10'sd494, 10'sd289, 12'sd1190}, {12'sd-1277, 11'sd-660, 7'sd-59}},
{{12'sd1327, 12'sd1697, 8'sd-67}, {10'sd372, 12'sd1802, 12'sd-1694}, {9'sd254, 11'sd-1009, 13'sd2611}},
{{12'sd-1279, 11'sd-855, 10'sd-319}, {13'sd-2786, 13'sd-2522, 11'sd827}, {14'sd-4328, 12'sd-1339, 12'sd1962}},
{{12'sd-1409, 10'sd-446, 11'sd919}, {11'sd970, 13'sd-2180, 13'sd2439}, {11'sd552, 12'sd-1130, 13'sd-2279}},
{{12'sd-1637, 11'sd-1011, 13'sd-2553}, {10'sd375, 12'sd-2014, 13'sd2449}, {12'sd1906, 12'sd1231, 11'sd785}},
{{12'sd-1157, 13'sd2107, 12'sd1460}, {12'sd1133, 11'sd-717, 13'sd2369}, {11'sd-936, 6'sd19, 13'sd2761}},
{{13'sd-3207, 13'sd-3548, 13'sd-2947}, {11'sd-910, 13'sd2522, 13'sd2436}, {10'sd439, 10'sd-394, 9'sd180}},
{{14'sd5455, 13'sd3191, 13'sd-2745}, {13'sd3243, 13'sd2397, 11'sd-762}, {12'sd1387, 7'sd38, 11'sd800}},
{{13'sd3226, 12'sd1626, 14'sd-5701}, {13'sd4064, 13'sd2716, 13'sd-2773}, {13'sd3598, 13'sd2075, 12'sd1360}},
{{11'sd-836, 12'sd-1577, 11'sd768}, {12'sd1278, 12'sd2029, 11'sd-857}, {12'sd-1495, 12'sd1337, 13'sd-2153}},
{{13'sd3490, 12'sd-1725, 8'sd-124}, {13'sd3603, 12'sd-1179, 11'sd837}, {10'sd379, 13'sd-3792, 13'sd-3449}},
{{12'sd-1076, 13'sd2278, 8'sd119}, {12'sd1913, 10'sd-282, 12'sd1032}, {13'sd-2204, 11'sd-637, 10'sd473}},
{{13'sd-2949, 10'sd456, 13'sd-2452}, {13'sd-2897, 12'sd-1690, 12'sd1940}, {13'sd3419, 12'sd-1993, 12'sd1644}},
{{12'sd-1508, 13'sd-2294, 13'sd2479}, {13'sd-3043, 13'sd-3163, 12'sd-1295}, {14'sd-5020, 13'sd-2426, 12'sd1222}}},
{
{{12'sd1711, 11'sd770, 13'sd3110}, {13'sd-2302, 11'sd-583, 13'sd2227}, {12'sd1956, 9'sd-175, 13'sd-3144}},
{{12'sd-2047, 13'sd2593, 11'sd654}, {8'sd-90, 13'sd-2163, 9'sd-249}, {11'sd-680, 13'sd2751, 13'sd2862}},
{{12'sd-2009, 11'sd-898, 12'sd-1834}, {10'sd337, 13'sd-3159, 5'sd8}, {13'sd-2790, 9'sd194, 11'sd696}},
{{13'sd2347, 12'sd-1307, 12'sd-1296}, {13'sd3329, 12'sd1152, 12'sd1974}, {13'sd-2356, 11'sd-934, 12'sd-1989}},
{{11'sd727, 11'sd-826, 11'sd871}, {12'sd-1151, 11'sd-995, 12'sd1561}, {12'sd-1261, 13'sd3055, 13'sd-3055}},
{{11'sd-915, 9'sd162, 13'sd4039}, {10'sd-397, 13'sd-2152, 13'sd3045}, {11'sd-786, 10'sd-323, 11'sd-840}},
{{14'sd-4362, 11'sd-766, 13'sd-3470}, {11'sd-589, 12'sd-1193, 13'sd-2394}, {13'sd3324, 14'sd5300, 12'sd1361}},
{{8'sd94, 12'sd1157, 12'sd2035}, {10'sd380, 13'sd2599, 10'sd-294}, {13'sd-3258, 13'sd2452, 12'sd1170}},
{{12'sd-1995, 11'sd-753, 13'sd2670}, {13'sd-2248, 11'sd-817, 13'sd2857}, {13'sd-2798, 6'sd-31, 12'sd1147}},
{{9'sd234, 8'sd85, 13'sd3328}, {11'sd851, 11'sd534, 12'sd1904}, {11'sd-839, 12'sd-1925, 11'sd-911}},
{{14'sd5675, 10'sd-277, 14'sd-5526}, {14'sd5071, 13'sd-2548, 14'sd-5856}, {12'sd-1421, 14'sd-4842, 13'sd-3602}},
{{11'sd608, 10'sd-268, 13'sd2328}, {13'sd-2779, 13'sd-2702, 13'sd2442}, {13'sd-3752, 12'sd1304, 11'sd567}},
{{13'sd-2451, 9'sd157, 13'sd2177}, {13'sd-3643, 10'sd489, 14'sd4985}, {13'sd-2339, 11'sd564, 13'sd3585}},
{{13'sd-2075, 8'sd109, 12'sd-1900}, {9'sd-166, 13'sd2249, 10'sd270}, {13'sd2098, 10'sd497, 11'sd717}},
{{10'sd453, 12'sd-1606, 12'sd1964}, {10'sd293, 8'sd99, 13'sd-2732}, {13'sd3493, 12'sd-1733, 13'sd2240}},
{{14'sd-4104, 10'sd402, 12'sd2009}, {13'sd-2961, 11'sd591, 13'sd3038}, {13'sd-3326, 11'sd-564, 13'sd3701}},
{{12'sd-1626, 13'sd2206, 12'sd1672}, {11'sd-808, 13'sd2468, 13'sd2387}, {10'sd417, 13'sd2473, 12'sd2031}},
{{14'sd-6536, 14'sd-5441, 13'sd2829}, {14'sd-5064, 11'sd882, 14'sd4971}, {13'sd3113, 13'sd3623, 14'sd4988}},
{{13'sd-3007, 12'sd1793, 11'sd-1013}, {6'sd-20, 12'sd1526, 10'sd-429}, {11'sd-658, 13'sd-2379, 13'sd2554}},
{{13'sd3949, 9'sd-143, 13'sd3932}, {10'sd338, 12'sd1368, 13'sd2496}, {10'sd-336, 11'sd893, 13'sd3071}},
{{11'sd792, 13'sd2896, 9'sd183}, {12'sd-1367, 12'sd1447, 12'sd-1298}, {12'sd1690, 12'sd1959, 12'sd1662}},
{{12'sd-1443, 11'sd864, 9'sd160}, {4'sd5, 10'sd414, 13'sd-3938}, {10'sd-429, 9'sd162, 13'sd-3811}},
{{12'sd-1628, 11'sd-693, 11'sd513}, {11'sd-637, 12'sd1155, 10'sd-508}, {13'sd2069, 12'sd-1200, 6'sd-20}},
{{12'sd-1717, 11'sd971, 12'sd1200}, {6'sd-24, 12'sd1965, 13'sd2084}, {11'sd-526, 11'sd1018, 11'sd-562}},
{{12'sd-1872, 13'sd2208, 13'sd2266}, {13'sd-2229, 12'sd-2018, 8'sd74}, {14'sd-5809, 13'sd-3994, 13'sd2053}},
{{13'sd-2178, 12'sd1947, 13'sd-2956}, {12'sd1193, 10'sd-400, 12'sd-1706}, {13'sd-2635, 12'sd1050, 13'sd2417}},
{{12'sd1806, 12'sd1948, 11'sd-820}, {8'sd-68, 10'sd-454, 11'sd861}, {9'sd135, 13'sd-2647, 12'sd1962}},
{{10'sd-308, 10'sd-303, 12'sd-1214}, {11'sd852, 13'sd3094, 11'sd-801}, {13'sd-2737, 12'sd1686, 10'sd423}},
{{12'sd-1948, 14'sd-4526, 14'sd-4433}, {11'sd567, 11'sd-820, 13'sd-3415}, {13'sd2167, 13'sd2304, 9'sd128}},
{{12'sd1323, 12'sd-1786, 12'sd1459}, {14'sd4453, 11'sd981, 7'sd39}, {13'sd2693, 11'sd-689, 9'sd230}},
{{12'sd-1087, 1'sd0, 13'sd2395}, {12'sd-1681, 13'sd-3364, 10'sd-405}, {11'sd-608, 8'sd-85, 12'sd1777}},
{{13'sd-2621, 13'sd-2273, 13'sd2744}, {10'sd-397, 9'sd-240, 12'sd-1475}, {11'sd749, 12'sd1798, 13'sd3568}},
{{9'sd-180, 13'sd2336, 11'sd943}, {12'sd1371, 11'sd-625, 12'sd1581}, {8'sd65, 8'sd-118, 13'sd-2144}},
{{13'sd3041, 5'sd15, 12'sd2022}, {13'sd-2654, 8'sd-100, 13'sd3250}, {11'sd714, 13'sd-2542, 11'sd-978}},
{{13'sd2497, 12'sd-1771, 11'sd688}, {10'sd-418, 13'sd-2516, 10'sd504}, {13'sd-3667, 12'sd-1223, 13'sd-2507}},
{{12'sd-1592, 12'sd-1751, 12'sd-1087}, {13'sd2177, 11'sd964, 12'sd1143}, {12'sd-1497, 11'sd836, 12'sd1593}},
{{12'sd-1876, 12'sd1375, 12'sd1544}, {12'sd1785, 12'sd1845, 9'sd228}, {11'sd928, 13'sd2156, 5'sd15}},
{{14'sd-4352, 11'sd556, 13'sd-2106}, {14'sd-4226, 7'sd-59, 12'sd-1211}, {12'sd1220, 13'sd3074, 12'sd1974}},
{{10'sd-328, 13'sd2077, 12'sd1855}, {11'sd-1012, 12'sd-1937, 13'sd-3365}, {13'sd3489, 13'sd2147, 11'sd-802}},
{{10'sd323, 11'sd-581, 13'sd-2698}, {10'sd321, 10'sd415, 12'sd-1663}, {11'sd532, 12'sd-1866, 12'sd1194}},
{{6'sd-29, 13'sd-2230, 13'sd2824}, {13'sd-2596, 10'sd471, 12'sd1815}, {12'sd1982, 13'sd2180, 12'sd1649}},
{{13'sd-3448, 11'sd807, 12'sd1947}, {10'sd284, 13'sd2497, 12'sd1715}, {13'sd-3356, 9'sd252, 8'sd89}},
{{12'sd1231, 12'sd1392, 8'sd-72}, {10'sd500, 11'sd953, 13'sd-3269}, {11'sd-768, 9'sd222, 13'sd2159}},
{{10'sd370, 8'sd-97, 13'sd2383}, {12'sd1257, 13'sd3583, 12'sd-1429}, {12'sd-1789, 10'sd-412, 8'sd-105}},
{{12'sd1900, 12'sd1107, 13'sd-2679}, {12'sd1588, 12'sd-1107, 11'sd767}, {12'sd1836, 11'sd526, 11'sd-646}},
{{11'sd-996, 13'sd2867, 13'sd2580}, {12'sd-1617, 11'sd945, 9'sd171}, {11'sd870, 9'sd168, 11'sd919}},
{{13'sd-2930, 13'sd-2618, 12'sd-1300}, {12'sd-1074, 11'sd-792, 12'sd-1634}, {14'sd4253, 11'sd792, 13'sd2512}},
{{11'sd-904, 12'sd-1616, 8'sd-110}, {12'sd-1051, 10'sd-310, 12'sd-1493}, {12'sd-1212, 12'sd-1203, 12'sd1162}},
{{13'sd-2099, 12'sd-1150, 10'sd-361}, {12'sd1728, 12'sd1558, 13'sd-2280}, {12'sd-1320, 13'sd-2348, 13'sd2125}},
{{11'sd897, 12'sd-1024, 12'sd1359}, {11'sd1014, 13'sd-2588, 13'sd-2364}, {11'sd772, 11'sd770, 12'sd-1050}},
{{13'sd2239, 13'sd-2269, 12'sd-1139}, {12'sd1217, 12'sd-1035, 13'sd2131}, {10'sd-311, 9'sd213, 11'sd-721}},
{{12'sd1596, 12'sd-1311, 12'sd1512}, {11'sd-745, 12'sd1847, 9'sd-192}, {11'sd-513, 11'sd857, 13'sd-3138}},
{{14'sd-5380, 14'sd-4393, 12'sd-1293}, {12'sd1609, 11'sd-720, 13'sd-3659}, {12'sd1483, 13'sd2177, 13'sd-2573}},
{{13'sd2084, 11'sd-593, 13'sd-2243}, {12'sd1840, 13'sd-2925, 12'sd-1980}, {12'sd-1303, 12'sd1517, 11'sd582}},
{{13'sd-2306, 11'sd886, 12'sd1875}, {12'sd-1249, 12'sd-1307, 13'sd-2466}, {13'sd2301, 11'sd903, 8'sd-127}},
{{11'sd-909, 11'sd995, 12'sd1515}, {11'sd529, 12'sd1322, 13'sd2496}, {12'sd1060, 10'sd271, 12'sd-1459}},
{{12'sd1853, 11'sd1021, 9'sd198}, {13'sd-3152, 12'sd-1483, 11'sd-750}, {13'sd-2683, 12'sd1313, 11'sd707}},
{{12'sd-2006, 12'sd-1060, 13'sd3207}, {13'sd-2614, 11'sd-987, 12'sd1884}, {9'sd-222, 14'sd4381, 14'sd5544}},
{{12'sd-1271, 13'sd-3341, 13'sd-3806}, {13'sd-2146, 13'sd2155, 13'sd-2202}, {10'sd-367, 13'sd2406, 10'sd333}},
{{13'sd-2613, 12'sd-1623, 13'sd-2182}, {12'sd-1738, 4'sd-7, 12'sd1551}, {12'sd1936, 12'sd-1138, 12'sd-1712}},
{{11'sd573, 9'sd-225, 9'sd181}, {13'sd-3361, 12'sd-1391, 13'sd2299}, {12'sd-1891, 8'sd102, 13'sd2573}},
{{9'sd-249, 12'sd-1256, 13'sd-2077}, {11'sd-959, 11'sd923, 13'sd2629}, {11'sd702, 12'sd1763, 11'sd853}},
{{8'sd-106, 12'sd-1411, 13'sd2855}, {12'sd1254, 12'sd1589, 13'sd3153}, {13'sd-2589, 5'sd11, 13'sd-2147}},
{{14'sd-4305, 8'sd-100, 13'sd-4058}, {13'sd2118, 13'sd3210, 11'sd-997}, {12'sd1423, 11'sd924, 13'sd-3158}}},
{
{{11'sd928, 11'sd-930, 12'sd-1287}, {10'sd320, 13'sd-2365, 11'sd912}, {10'sd-332, 12'sd-1273, 4'sd7}},
{{12'sd1564, 11'sd-938, 12'sd1738}, {12'sd-2012, 10'sd-291, 12'sd-1782}, {12'sd-1151, 12'sd-1932, 13'sd-2421}},
{{10'sd-457, 11'sd916, 10'sd-437}, {13'sd2205, 9'sd-155, 10'sd-278}, {12'sd-1249, 13'sd-3327, 13'sd-2248}},
{{12'sd1965, 11'sd548, 13'sd2240}, {12'sd1446, 12'sd1213, 13'sd2086}, {12'sd1648, 10'sd-387, 12'sd1286}},
{{9'sd223, 10'sd-435, 13'sd2524}, {12'sd-1562, 13'sd-2296, 13'sd2275}, {12'sd1462, 12'sd-1610, 12'sd1427}},
{{10'sd-317, 12'sd-1309, 12'sd1461}, {13'sd2102, 11'sd573, 12'sd-1956}, {8'sd93, 13'sd3016, 11'sd-795}},
{{13'sd2660, 13'sd-2397, 13'sd-2551}, {12'sd1204, 11'sd-597, 11'sd626}, {12'sd1291, 13'sd-2121, 12'sd1523}},
{{10'sd394, 11'sd-822, 13'sd2749}, {11'sd-842, 12'sd1931, 10'sd291}, {12'sd-1078, 12'sd-1288, 13'sd-2164}},
{{12'sd1218, 13'sd2090, 13'sd-2515}, {12'sd-1689, 13'sd2103, 11'sd769}, {7'sd58, 12'sd1370, 12'sd-1439}},
{{12'sd-1784, 12'sd-1897, 13'sd-2875}, {13'sd-2616, 13'sd-2299, 8'sd126}, {13'sd-2164, 8'sd89, 12'sd-1333}},
{{12'sd1876, 12'sd1324, 11'sd-757}, {12'sd1801, 13'sd3776, 13'sd3405}, {13'sd2123, 13'sd2391, 13'sd2205}},
{{12'sd1544, 12'sd1279, 13'sd2227}, {12'sd1538, 13'sd-2503, 12'sd-1334}, {12'sd1929, 12'sd1168, 13'sd2187}},
{{10'sd-378, 11'sd-623, 13'sd-2215}, {11'sd-961, 13'sd-2745, 10'sd458}, {11'sd-973, 12'sd1874, 12'sd-1297}},
{{11'sd864, 11'sd916, 10'sd-412}, {13'sd-2405, 11'sd-1003, 10'sd337}, {10'sd-298, 13'sd2073, 12'sd-1983}},
{{12'sd1802, 13'sd2351, 11'sd-959}, {10'sd287, 13'sd-2621, 12'sd-1612}, {12'sd1111, 10'sd363, 11'sd840}},
{{13'sd2533, 10'sd291, 12'sd1697}, {13'sd-2519, 12'sd-1543, 12'sd-1414}, {13'sd2397, 10'sd-511, 13'sd2573}},
{{12'sd-1629, 11'sd-993, 12'sd-1051}, {11'sd-799, 12'sd-1693, 12'sd1190}, {11'sd652, 7'sd-50, 13'sd-2655}},
{{13'sd2107, 13'sd3418, 13'sd-2731}, {12'sd1448, 13'sd-3057, 13'sd-3368}, {12'sd-1293, 9'sd-194, 13'sd-4064}},
{{12'sd-1216, 9'sd-238, 11'sd-746}, {12'sd-1814, 10'sd-480, 11'sd552}, {9'sd177, 11'sd548, 12'sd-1856}},
{{12'sd-1308, 10'sd378, 11'sd-528}, {10'sd510, 13'sd-2610, 13'sd-2692}, {12'sd1344, 12'sd1540, 11'sd817}},
{{10'sd347, 13'sd-2833, 12'sd-1962}, {12'sd-1392, 7'sd-38, 11'sd906}, {12'sd-1965, 12'sd1197, 12'sd1186}},
{{12'sd-1741, 11'sd-763, 11'sd-838}, {13'sd-2740, 13'sd-2093, 12'sd1264}, {13'sd2633, 11'sd-679, 12'sd-1290}},
{{11'sd-611, 12'sd1605, 12'sd-1922}, {12'sd1147, 13'sd2276, 12'sd-1640}, {12'sd-1683, 10'sd315, 12'sd1113}},
{{12'sd1908, 11'sd729, 11'sd975}, {13'sd2516, 11'sd754, 13'sd2457}, {10'sd327, 13'sd2681, 12'sd-1052}},
{{13'sd-2964, 10'sd504, 13'sd-2409}, {13'sd2317, 13'sd2392, 12'sd1267}, {12'sd-1833, 11'sd-863, 11'sd-809}},
{{12'sd-1550, 12'sd1635, 13'sd2512}, {9'sd-234, 12'sd1717, 12'sd1767}, {12'sd1872, 12'sd-1538, 12'sd1250}},
{{7'sd38, 13'sd2544, 9'sd-184}, {13'sd2720, 11'sd576, 12'sd1690}, {12'sd1985, 11'sd532, 12'sd1342}},
{{13'sd-2267, 13'sd2842, 13'sd-3016}, {10'sd-266, 13'sd-2297, 12'sd-1671}, {8'sd-111, 12'sd-1045, 12'sd-1185}},
{{11'sd-684, 13'sd2568, 13'sd2132}, {13'sd-2516, 9'sd-164, 13'sd-2129}, {11'sd938, 10'sd498, 9'sd202}},
{{6'sd-21, 13'sd-3052, 10'sd-261}, {11'sd880, 12'sd1632, 10'sd-261}, {11'sd907, 12'sd1518, 12'sd-1109}},
{{11'sd925, 11'sd-803, 12'sd-1878}, {10'sd322, 12'sd-1738, 11'sd-762}, {13'sd-2497, 12'sd-1737, 13'sd-2517}},
{{11'sd881, 12'sd-1211, 12'sd1949}, {12'sd1396, 11'sd655, 12'sd1663}, {12'sd1051, 10'sd304, 12'sd-1553}},
{{12'sd1195, 12'sd-1434, 12'sd-1616}, {13'sd2824, 11'sd-675, 11'sd585}, {8'sd94, 12'sd1682, 12'sd-1510}},
{{8'sd88, 13'sd2244, 13'sd2417}, {10'sd472, 12'sd1303, 12'sd-1903}, {13'sd-2566, 11'sd743, 5'sd-12}},
{{10'sd-464, 12'sd-1625, 13'sd-2207}, {10'sd357, 11'sd659, 11'sd-833}, {12'sd-1195, 12'sd-1318, 13'sd2827}},
{{12'sd1256, 12'sd-1893, 9'sd242}, {10'sd310, 11'sd-909, 12'sd-1348}, {11'sd529, 12'sd1471, 10'sd-291}},
{{12'sd1392, 9'sd-242, 12'sd1136}, {10'sd-324, 10'sd-423, 11'sd-729}, {8'sd-100, 10'sd436, 12'sd-1805}},
{{11'sd-933, 12'sd-1242, 12'sd-1270}, {11'sd-1018, 12'sd1388, 13'sd-2589}, {12'sd2005, 9'sd206, 12'sd1097}},
{{13'sd2133, 12'sd2033, 13'sd-2812}, {12'sd1702, 12'sd1923, 13'sd-2143}, {10'sd299, 13'sd2630, 8'sd114}},
{{13'sd2252, 12'sd1223, 12'sd1042}, {12'sd1781, 8'sd-115, 11'sd-665}, {11'sd-878, 10'sd337, 11'sd-898}},
{{10'sd381, 8'sd104, 12'sd1785}, {12'sd1602, 12'sd-1247, 12'sd-1697}, {12'sd-2025, 11'sd-753, 12'sd-1586}},
{{12'sd-1478, 13'sd2066, 10'sd-362}, {13'sd2558, 11'sd591, 12'sd-1154}, {11'sd884, 10'sd309, 12'sd1448}},
{{12'sd-1341, 12'sd1391, 12'sd1552}, {12'sd1671, 12'sd1381, 13'sd2541}, {12'sd1275, 9'sd-226, 12'sd-1063}},
{{12'sd-2019, 12'sd-1935, 12'sd-1848}, {13'sd2163, 12'sd1277, 12'sd1863}, {12'sd-1396, 12'sd-1743, 10'sd-497}},
{{11'sd-757, 10'sd-468, 11'sd958}, {12'sd1372, 12'sd2043, 8'sd-124}, {12'sd1426, 11'sd958, 12'sd-1704}},
{{13'sd2409, 11'sd735, 12'sd-1362}, {10'sd-298, 11'sd783, 10'sd386}, {6'sd-26, 11'sd721, 12'sd-1951}},
{{10'sd508, 11'sd-583, 8'sd-81}, {13'sd-2426, 11'sd-803, 12'sd1113}, {10'sd257, 10'sd-398, 13'sd-2321}},
{{12'sd-1106, 12'sd1600, 12'sd-1889}, {11'sd666, 10'sd502, 12'sd1723}, {13'sd-2551, 12'sd-1356, 13'sd-2906}},
{{12'sd1810, 13'sd-2330, 13'sd2115}, {13'sd-2336, 9'sd-214, 11'sd-548}, {12'sd1415, 11'sd999, 10'sd447}},
{{13'sd-2604, 11'sd-586, 12'sd1198}, {12'sd-1827, 12'sd1141, 11'sd-847}, {13'sd-2623, 13'sd2245, 12'sd1602}},
{{11'sd823, 11'sd920, 12'sd1641}, {12'sd-1194, 10'sd459, 12'sd-1464}, {8'sd124, 12'sd1650, 10'sd-280}},
{{11'sd823, 12'sd-1947, 12'sd1774}, {9'sd-224, 12'sd1249, 12'sd1563}, {12'sd-1971, 12'sd1396, 11'sd515}},
{{12'sd-2011, 13'sd-2551, 11'sd694}, {12'sd2000, 11'sd-570, 12'sd-1189}, {12'sd1647, 12'sd1119, 13'sd-2572}},
{{13'sd2096, 11'sd-539, 10'sd413}, {10'sd476, 13'sd2256, 13'sd-2736}, {12'sd-2019, 13'sd-2212, 10'sd-476}},
{{9'sd-156, 13'sd2309, 12'sd-1376}, {13'sd2391, 13'sd2559, 12'sd-1473}, {12'sd2030, 9'sd157, 11'sd687}},
{{6'sd-24, 11'sd-888, 9'sd-205}, {13'sd-2476, 13'sd2810, 11'sd658}, {11'sd763, 11'sd-513, 12'sd1074}},
{{8'sd91, 13'sd3122, 13'sd-2061}, {12'sd-1599, 12'sd1493, 13'sd-2254}, {11'sd722, 11'sd866, 11'sd-765}},
{{13'sd2077, 12'sd1783, 11'sd951}, {13'sd2567, 11'sd-651, 13'sd-2294}, {7'sd36, 12'sd-1331, 11'sd-759}},
{{12'sd1377, 7'sd54, 12'sd1367}, {8'sd-111, 11'sd-847, 13'sd2981}, {13'sd2418, 9'sd170, 13'sd2875}},
{{12'sd1086, 12'sd1604, 13'sd-2323}, {13'sd2641, 13'sd-2059, 13'sd-2782}, {12'sd-1857, 12'sd1277, 11'sd-861}},
{{12'sd1946, 11'sd905, 9'sd202}, {11'sd944, 13'sd-2689, 11'sd-635}, {12'sd-1130, 13'sd2797, 13'sd-2166}},
{{12'sd1152, 11'sd-682, 10'sd-357}, {13'sd2050, 11'sd-911, 11'sd-879}, {12'sd-2039, 10'sd-259, 12'sd-1534}},
{{11'sd716, 10'sd267, 12'sd-1741}, {13'sd2628, 3'sd3, 13'sd2306}, {11'sd-980, 13'sd-2505, 13'sd-2800}},
{{13'sd2488, 13'sd2303, 12'sd-1066}, {11'sd654, 13'sd-2405, 13'sd2109}, {10'sd-305, 13'sd-2543, 7'sd-48}}},
{
{{13'sd2437, 12'sd-1407, 11'sd736}, {12'sd-1529, 12'sd1508, 12'sd1397}, {12'sd-1886, 10'sd-433, 11'sd793}},
{{13'sd-3119, 10'sd499, 11'sd-553}, {12'sd-1522, 12'sd-1954, 13'sd-2493}, {9'sd180, 13'sd2425, 12'sd1242}},
{{13'sd-2090, 13'sd2350, 12'sd1024}, {12'sd-1286, 13'sd2561, 12'sd-1844}, {10'sd-499, 12'sd1083, 11'sd548}},
{{11'sd558, 12'sd1664, 11'sd-1018}, {12'sd-1965, 13'sd2690, 13'sd-2178}, {12'sd-1962, 12'sd-1547, 9'sd-242}},
{{11'sd-763, 12'sd1495, 12'sd-1312}, {11'sd-646, 11'sd-514, 11'sd-1011}, {11'sd-552, 12'sd-1027, 11'sd-601}},
{{11'sd-797, 12'sd1910, 11'sd637}, {10'sd-375, 13'sd-2374, 5'sd-12}, {12'sd1623, 7'sd52, 12'sd2043}},
{{12'sd1497, 11'sd772, 11'sd-931}, {9'sd248, 7'sd60, 11'sd-829}, {13'sd2491, 12'sd1289, 8'sd86}},
{{12'sd-1555, 13'sd3143, 12'sd1081}, {13'sd2175, 13'sd2592, 12'sd1694}, {13'sd-2494, 13'sd-2330, 12'sd1495}},
{{6'sd20, 12'sd-1574, 10'sd499}, {12'sd-1734, 10'sd385, 12'sd-1259}, {12'sd-1224, 11'sd841, 13'sd2949}},
{{11'sd844, 10'sd280, 10'sd322}, {10'sd304, 11'sd-743, 12'sd1798}, {12'sd-1485, 10'sd481, 13'sd-2281}},
{{14'sd5085, 12'sd1968, 13'sd-2957}, {12'sd1759, 8'sd71, 11'sd-937}, {13'sd3456, 10'sd-488, 12'sd1352}},
{{11'sd-798, 12'sd-1728, 8'sd-97}, {12'sd1578, 10'sd439, 12'sd-1853}, {11'sd1022, 13'sd-2166, 9'sd-142}},
{{13'sd2497, 13'sd-2704, 12'sd-1486}, {12'sd1067, 12'sd-1727, 12'sd1906}, {12'sd1900, 12'sd-1130, 12'sd-1184}},
{{13'sd2479, 12'sd1578, 13'sd-2123}, {8'sd-122, 13'sd-2126, 6'sd25}, {13'sd-2708, 12'sd-1305, 13'sd-2755}},
{{12'sd-1487, 12'sd-1215, 10'sd-506}, {12'sd-1607, 11'sd-789, 11'sd-908}, {11'sd979, 12'sd-1805, 12'sd1120}},
{{12'sd-1359, 9'sd-227, 11'sd-903}, {12'sd1808, 12'sd-1247, 13'sd-2235}, {12'sd-1298, 13'sd2213, 10'sd-460}},
{{13'sd-2314, 12'sd1082, 11'sd535}, {12'sd-1698, 11'sd716, 5'sd8}, {12'sd-1962, 11'sd-896, 11'sd960}},
{{13'sd-3276, 13'sd-2426, 6'sd-29}, {11'sd908, 13'sd-2749, 13'sd3426}, {13'sd3057, 13'sd2438, 11'sd832}},
{{11'sd-676, 8'sd-81, 13'sd-2731}, {11'sd976, 13'sd-2260, 12'sd-1468}, {8'sd-91, 13'sd2532, 12'sd-1770}},
{{11'sd572, 13'sd-2370, 11'sd867}, {11'sd743, 10'sd-276, 12'sd-1247}, {12'sd-1596, 11'sd-1001, 13'sd-2723}},
{{11'sd528, 10'sd433, 11'sd-737}, {12'sd1375, 13'sd-2103, 11'sd-830}, {13'sd2075, 13'sd2151, 11'sd881}},
{{13'sd-2391, 13'sd-2335, 12'sd-1991}, {8'sd-85, 11'sd-951, 12'sd-1730}, {9'sd-141, 11'sd620, 11'sd-713}},
{{12'sd-1540, 11'sd-619, 11'sd-974}, {12'sd1752, 13'sd2121, 11'sd-725}, {9'sd195, 13'sd-2892, 12'sd-1873}},
{{11'sd694, 9'sd212, 9'sd247}, {10'sd278, 12'sd-1370, 12'sd-1759}, {12'sd-1767, 12'sd-1854, 9'sd-234}},
{{11'sd-546, 12'sd-2016, 11'sd889}, {13'sd-3014, 13'sd2053, 13'sd3418}, {11'sd946, 11'sd541, 12'sd1183}},
{{13'sd3111, 11'sd-587, 12'sd1622}, {12'sd1446, 11'sd793, 12'sd1075}, {10'sd-272, 11'sd-707, 12'sd1909}},
{{13'sd-2222, 11'sd-777, 13'sd-2810}, {12'sd1634, 13'sd2891, 9'sd253}, {13'sd2387, 13'sd2818, 11'sd1005}},
{{13'sd2375, 12'sd-1437, 11'sd559}, {8'sd-105, 8'sd114, 12'sd2025}, {11'sd-589, 12'sd1206, 12'sd-1492}},
{{11'sd795, 13'sd-2472, 12'sd-1686}, {12'sd1270, 12'sd-1282, 13'sd-2650}, {11'sd562, 9'sd166, 12'sd1331}},
{{11'sd-592, 12'sd-1191, 11'sd-809}, {12'sd1880, 12'sd1867, 11'sd-970}, {13'sd-3493, 12'sd-1482, 11'sd655}},
{{13'sd2486, 13'sd2069, 3'sd-3}, {11'sd1004, 11'sd-648, 13'sd2184}, {13'sd-2715, 13'sd-2640, 11'sd709}},
{{13'sd2195, 13'sd-2054, 11'sd967}, {3'sd2, 12'sd-1945, 12'sd-1078}, {12'sd-1194, 11'sd631, 11'sd525}},
{{12'sd1173, 13'sd2147, 9'sd-171}, {12'sd-1190, 10'sd-439, 12'sd1756}, {12'sd-1869, 10'sd-450, 11'sd770}},
{{12'sd2005, 9'sd186, 10'sd308}, {11'sd886, 11'sd610, 6'sd17}, {8'sd-113, 13'sd2621, 12'sd1896}},
{{10'sd468, 12'sd1819, 9'sd138}, {7'sd-60, 12'sd1154, 8'sd-91}, {10'sd-356, 13'sd-2193, 11'sd-1014}},
{{12'sd1181, 13'sd2590, 13'sd2556}, {11'sd887, 6'sd31, 12'sd-1915}, {13'sd2516, 12'sd-1185, 12'sd1978}},
{{13'sd2661, 11'sd-551, 10'sd-285}, {8'sd-95, 12'sd-1321, 12'sd-2033}, {9'sd-203, 9'sd193, 12'sd-1336}},
{{1'sd0, 12'sd-1991, 11'sd-987}, {13'sd-3465, 9'sd255, 13'sd-3378}, {13'sd-2436, 9'sd185, 11'sd-770}},
{{12'sd-1837, 13'sd-2255, 8'sd97}, {9'sd-202, 12'sd1453, 11'sd955}, {12'sd1433, 11'sd-917, 7'sd38}},
{{13'sd2415, 13'sd2513, 13'sd2269}, {12'sd-1317, 12'sd-1350, 13'sd-2751}, {11'sd-776, 12'sd-1913, 13'sd2906}},
{{13'sd-2834, 12'sd1759, 11'sd-863}, {12'sd-2043, 12'sd1104, 13'sd-2534}, {12'sd-1131, 13'sd2314, 12'sd1288}},
{{11'sd-742, 12'sd-1812, 11'sd597}, {11'sd740, 12'sd-1239, 13'sd2262}, {13'sd-2410, 11'sd-585, 12'sd1274}},
{{11'sd-605, 10'sd292, 11'sd992}, {12'sd-1716, 12'sd-1787, 11'sd904}, {12'sd-1719, 11'sd567, 12'sd-1459}},
{{10'sd387, 10'sd510, 12'sd1285}, {11'sd580, 11'sd-904, 12'sd1064}, {13'sd2632, 13'sd-2265, 12'sd-1348}},
{{12'sd1980, 12'sd1796, 12'sd-1905}, {12'sd-1694, 9'sd-179, 13'sd2097}, {12'sd1840, 11'sd742, 12'sd-1561}},
{{12'sd1192, 13'sd-2583, 10'sd-322}, {11'sd634, 11'sd657, 12'sd-1158}, {12'sd2016, 11'sd549, 9'sd-196}},
{{13'sd2137, 13'sd2742, 12'sd-1270}, {7'sd45, 13'sd2620, 13'sd-2093}, {7'sd53, 13'sd2756, 12'sd1947}},
{{13'sd-2615, 8'sd-65, 10'sd372}, {11'sd-578, 10'sd-367, 11'sd957}, {12'sd1781, 13'sd-2745, 12'sd-1611}},
{{10'sd-501, 11'sd808, 13'sd-2939}, {12'sd-1199, 12'sd-1577, 12'sd1588}, {12'sd1378, 10'sd-410, 10'sd391}},
{{13'sd-2465, 12'sd1041, 13'sd2372}, {13'sd-2588, 11'sd877, 12'sd-1908}, {12'sd1522, 12'sd-1901, 11'sd872}},
{{13'sd2550, 9'sd-192, 12'sd1879}, {8'sd-115, 13'sd2338, 12'sd-1091}, {11'sd639, 12'sd-1314, 12'sd1601}},
{{12'sd1217, 11'sd-1000, 12'sd1843}, {11'sd720, 12'sd-1375, 12'sd1484}, {12'sd-2027, 10'sd339, 9'sd131}},
{{11'sd600, 12'sd1852, 11'sd604}, {12'sd-1566, 13'sd-2162, 12'sd-1457}, {12'sd1927, 13'sd2825, 13'sd3094}},
{{13'sd-2799, 12'sd-1642, 10'sd-392}, {11'sd-936, 13'sd2214, 13'sd-2625}, {12'sd-1366, 13'sd-2190, 12'sd2001}},
{{12'sd1840, 10'sd-504, 12'sd-1133}, {12'sd-1032, 11'sd-833, 10'sd-270}, {13'sd-3070, 11'sd758, 12'sd-1338}},
{{11'sd-578, 13'sd-2731, 9'sd-133}, {10'sd505, 12'sd-1024, 9'sd144}, {12'sd-1759, 7'sd55, 8'sd-73}},
{{12'sd1867, 11'sd884, 12'sd-1352}, {12'sd-2016, 10'sd330, 12'sd1884}, {12'sd1890, 11'sd-866, 13'sd2708}},
{{13'sd2104, 10'sd399, 12'sd-1174}, {12'sd1768, 12'sd1483, 11'sd-983}, {12'sd1147, 7'sd43, 13'sd3601}},
{{13'sd2218, 11'sd-969, 10'sd497}, {11'sd592, 12'sd1848, 11'sd981}, {10'sd346, 12'sd-1644, 11'sd-557}},
{{11'sd1016, 13'sd2651, 12'sd1165}, {11'sd783, 13'sd2394, 12'sd1203}, {13'sd2613, 12'sd1236, 10'sd-291}},
{{12'sd-1781, 13'sd2367, 3'sd3}, {11'sd730, 11'sd857, 8'sd-106}, {13'sd-3052, 12'sd-1032, 12'sd-1330}},
{{13'sd2770, 11'sd-732, 5'sd10}, {13'sd-2408, 12'sd-1240, 11'sd-783}, {11'sd862, 12'sd1061, 11'sd756}},
{{13'sd-2232, 12'sd-1772, 11'sd881}, {10'sd297, 11'sd-648, 12'sd-1865}, {10'sd-369, 13'sd-2139, 11'sd681}},
{{13'sd-2865, 12'sd-1315, 12'sd-1374}, {11'sd-531, 11'sd-865, 13'sd-2706}, {10'sd321, 10'sd256, 12'sd1428}}},
{
{{11'sd812, 12'sd-1759, 11'sd-856}, {10'sd-358, 12'sd-1199, 12'sd1162}, {11'sd956, 13'sd2294, 13'sd-2343}},
{{13'sd2320, 12'sd2001, 12'sd1618}, {12'sd1674, 12'sd-1093, 13'sd-2397}, {11'sd-513, 12'sd1791, 13'sd2483}},
{{12'sd1162, 10'sd491, 12'sd1376}, {12'sd-1097, 12'sd1609, 13'sd-2280}, {12'sd-1392, 12'sd-1494, 13'sd-3951}},
{{12'sd-1506, 13'sd-2785, 11'sd707}, {13'sd-2586, 13'sd-2075, 11'sd1011}, {11'sd592, 8'sd66, 11'sd-911}},
{{10'sd270, 13'sd-2873, 13'sd2466}, {13'sd2964, 13'sd2225, 13'sd2070}, {13'sd2650, 12'sd1188, 7'sd52}},
{{12'sd1758, 12'sd1349, 11'sd-624}, {11'sd-697, 12'sd-1184, 9'sd232}, {6'sd21, 10'sd259, 10'sd-408}},
{{10'sd-448, 11'sd797, 13'sd-2343}, {12'sd1163, 12'sd-1224, 13'sd2196}, {12'sd-1512, 13'sd-2091, 12'sd-1966}},
{{11'sd-949, 11'sd573, 12'sd1279}, {13'sd2325, 10'sd-323, 12'sd1790}, {13'sd3328, 12'sd1457, 12'sd-1721}},
{{13'sd-2489, 11'sd-915, 13'sd2141}, {12'sd-1929, 10'sd-332, 10'sd-428}, {12'sd1042, 11'sd-794, 9'sd-254}},
{{12'sd1338, 11'sd530, 12'sd-1138}, {12'sd-1641, 10'sd-395, 12'sd1695}, {12'sd1574, 13'sd-2237, 12'sd1932}},
{{12'sd-1601, 12'sd1554, 10'sd283}, {8'sd103, 10'sd-297, 13'sd3543}, {13'sd3302, 12'sd-1070, 13'sd2870}},
{{12'sd1617, 13'sd-2412, 10'sd436}, {13'sd2557, 12'sd-1542, 13'sd-2509}, {12'sd1103, 12'sd-1753, 8'sd-124}},
{{12'sd-1643, 9'sd-148, 12'sd-1654}, {12'sd-1886, 12'sd1270, 13'sd-2976}, {10'sd329, 11'sd906, 12'sd1367}},
{{12'sd1922, 12'sd-1945, 12'sd1583}, {9'sd-202, 13'sd2059, 12'sd1117}, {12'sd1318, 11'sd-720, 11'sd660}},
{{13'sd-2521, 11'sd944, 11'sd-822}, {12'sd1505, 12'sd1420, 9'sd231}, {12'sd1973, 12'sd-2002, 12'sd-1438}},
{{12'sd-1357, 12'sd-1161, 10'sd450}, {11'sd-639, 11'sd643, 9'sd171}, {11'sd-935, 11'sd908, 12'sd-1376}},
{{11'sd-637, 11'sd570, 11'sd-634}, {12'sd-1173, 13'sd2798, 11'sd-616}, {11'sd-960, 13'sd-2239, 11'sd-665}},
{{13'sd3853, 10'sd-505, 11'sd-1010}, {11'sd520, 11'sd-595, 11'sd-544}, {9'sd-201, 13'sd-3007, 13'sd-2409}},
{{11'sd-857, 9'sd-226, 12'sd-1484}, {13'sd2747, 11'sd-640, 7'sd48}, {12'sd1128, 12'sd-1618, 13'sd-2773}},
{{12'sd1242, 10'sd-441, 13'sd2889}, {13'sd2744, 12'sd-1183, 13'sd-2161}, {13'sd2321, 13'sd2055, 11'sd-685}},
{{8'sd113, 12'sd1939, 10'sd-322}, {12'sd-1740, 13'sd-2264, 5'sd12}, {12'sd-1960, 13'sd-2655, 13'sd2510}},
{{11'sd-775, 13'sd2398, 11'sd-569}, {10'sd-397, 11'sd-740, 10'sd335}, {13'sd2053, 12'sd1942, 11'sd941}},
{{13'sd2429, 13'sd-2134, 12'sd1750}, {12'sd-1875, 12'sd-1159, 13'sd-2548}, {10'sd-278, 12'sd1764, 8'sd-64}},
{{9'sd-231, 10'sd459, 11'sd-686}, {7'sd38, 13'sd-2358, 11'sd-713}, {12'sd-1501, 11'sd-1019, 11'sd679}},
{{11'sd-886, 11'sd-854, 12'sd-1586}, {12'sd-1937, 12'sd1622, 11'sd515}, {11'sd-885, 13'sd-3076, 11'sd-818}},
{{12'sd-2018, 12'sd1212, 11'sd667}, {13'sd2752, 12'sd-1071, 13'sd2538}, {12'sd-1192, 11'sd607, 12'sd-1444}},
{{11'sd698, 13'sd-2200, 9'sd204}, {12'sd-2019, 13'sd-2450, 12'sd-1338}, {12'sd-1369, 13'sd-2615, 10'sd386}},
{{10'sd-363, 11'sd-605, 12'sd-1517}, {13'sd-2326, 12'sd-1054, 13'sd-2719}, {12'sd2012, 6'sd-31, 11'sd900}},
{{11'sd663, 13'sd-2539, 13'sd2511}, {11'sd-787, 12'sd-1970, 11'sd-512}, {13'sd-2320, 11'sd663, 13'sd2969}},
{{9'sd-219, 13'sd2085, 12'sd1948}, {10'sd-424, 13'sd3043, 11'sd969}, {11'sd-872, 13'sd3307, 12'sd1931}},
{{12'sd1694, 10'sd441, 11'sd929}, {11'sd-659, 6'sd-31, 13'sd2173}, {13'sd2596, 12'sd-1462, 13'sd2125}},
{{11'sd888, 12'sd-1242, 10'sd-441}, {10'sd399, 12'sd1969, 13'sd-2898}, {13'sd-3198, 13'sd-2488, 13'sd-2087}},
{{10'sd-300, 13'sd-2573, 2'sd-1}, {13'sd2101, 13'sd2585, 13'sd-2355}, {10'sd278, 13'sd2172, 13'sd-2947}},
{{12'sd-1609, 11'sd732, 13'sd2213}, {11'sd-615, 9'sd-205, 13'sd2455}, {12'sd-1401, 10'sd337, 9'sd-196}},
{{12'sd1682, 8'sd-100, 12'sd-1203}, {9'sd-251, 13'sd-2233, 10'sd-422}, {12'sd1027, 13'sd-2229, 11'sd982}},
{{9'sd129, 10'sd-505, 12'sd-1516}, {12'sd1245, 12'sd2012, 12'sd1300}, {13'sd2703, 13'sd2462, 12'sd-1839}},
{{13'sd2426, 13'sd-2549, 10'sd-261}, {13'sd2408, 9'sd190, 12'sd1926}, {9'sd-171, 7'sd-35, 12'sd-1473}},
{{11'sd571, 13'sd-2429, 12'sd-1816}, {9'sd244, 13'sd-3091, 11'sd-797}, {12'sd1853, 13'sd-2730, 13'sd-2755}},
{{12'sd1586, 11'sd899, 13'sd3201}, {11'sd925, 12'sd1246, 13'sd3054}, {10'sd448, 10'sd358, 12'sd1802}},
{{13'sd-2406, 11'sd650, 13'sd-2145}, {11'sd-838, 12'sd1492, 13'sd-2427}, {13'sd2380, 13'sd2304, 8'sd-124}},
{{10'sd335, 12'sd2012, 13'sd2449}, {13'sd2174, 11'sd-800, 9'sd151}, {12'sd-1418, 9'sd-211, 12'sd-1683}},
{{11'sd708, 12'sd-1874, 13'sd-2460}, {13'sd2469, 7'sd55, 12'sd1675}, {11'sd-813, 9'sd-197, 12'sd-1309}},
{{12'sd1480, 12'sd-2038, 13'sd-2211}, {12'sd-1344, 12'sd-1459, 7'sd-40}, {13'sd2663, 12'sd-1661, 12'sd-1177}},
{{13'sd2770, 13'sd-2126, 13'sd-2666}, {12'sd1422, 12'sd1072, 11'sd-682}, {13'sd2747, 13'sd3922, 11'sd609}},
{{11'sd914, 12'sd1846, 12'sd1556}, {12'sd-1126, 10'sd-445, 11'sd762}, {12'sd1946, 13'sd-2283, 11'sd567}},
{{12'sd-1181, 12'sd1948, 12'sd1625}, {12'sd-1593, 12'sd-1171, 11'sd-898}, {13'sd-2373, 13'sd-2799, 13'sd-2763}},
{{11'sd808, 13'sd2053, 12'sd-2010}, {12'sd-1393, 12'sd-1576, 12'sd1642}, {13'sd-3097, 11'sd-993, 9'sd-158}},
{{10'sd489, 13'sd2510, 13'sd2455}, {12'sd-1354, 11'sd-853, 10'sd-310}, {12'sd-1243, 12'sd1347, 10'sd-373}},
{{11'sd680, 12'sd2028, 10'sd-307}, {12'sd1533, 12'sd1422, 11'sd-996}, {13'sd-2215, 12'sd1960, 11'sd-993}},
{{13'sd-2661, 12'sd1423, 12'sd1697}, {13'sd-2495, 12'sd1744, 13'sd-2357}, {12'sd1463, 11'sd891, 12'sd-1384}},
{{12'sd-2032, 11'sd-917, 10'sd-343}, {12'sd2047, 12'sd1936, 9'sd-165}, {12'sd1921, 12'sd1928, 12'sd1842}},
{{13'sd2872, 12'sd1806, 11'sd-695}, {12'sd-2014, 12'sd1983, 11'sd-631}, {12'sd1930, 12'sd-1212, 11'sd-631}},
{{12'sd-1480, 7'sd-58, 12'sd1209}, {12'sd1688, 13'sd-2710, 12'sd1186}, {12'sd-1916, 14'sd-4325, 12'sd-1640}},
{{11'sd526, 12'sd-1326, 11'sd851}, {12'sd1629, 13'sd-2345, 12'sd2020}, {10'sd-459, 11'sd989, 11'sd-582}},
{{11'sd917, 10'sd-452, 13'sd-2063}, {11'sd530, 13'sd-2389, 8'sd125}, {10'sd307, 11'sd893, 12'sd-1831}},
{{12'sd1715, 13'sd-2597, 12'sd1943}, {12'sd-1617, 11'sd-1012, 12'sd1615}, {13'sd2153, 9'sd-144, 13'sd2264}},
{{12'sd-1725, 12'sd-1749, 10'sd282}, {9'sd199, 12'sd1835, 13'sd-2330}, {11'sd-988, 13'sd2276, 6'sd-19}},
{{12'sd-1875, 13'sd2510, 10'sd491}, {13'sd-2323, 11'sd582, 12'sd1488}, {13'sd-2576, 2'sd1, 12'sd-1823}},
{{11'sd669, 13'sd-3067, 9'sd-169}, {13'sd2183, 12'sd-1051, 13'sd-3940}, {13'sd2715, 13'sd2436, 13'sd-2396}},
{{11'sd-942, 13'sd2585, 12'sd-1565}, {10'sd488, 13'sd2211, 13'sd2307}, {9'sd-255, 10'sd-379, 12'sd-1421}},
{{13'sd2517, 12'sd1704, 12'sd1148}, {11'sd629, 12'sd1859, 12'sd-1444}, {12'sd1726, 12'sd-1407, 11'sd911}},
{{13'sd2414, 13'sd2349, 12'sd-1342}, {13'sd-2135, 12'sd1957, 12'sd-1175}, {11'sd-546, 12'sd-1866, 12'sd-1885}},
{{12'sd-1849, 12'sd1495, 11'sd890}, {11'sd-657, 12'sd1430, 12'sd1787}, {13'sd2093, 11'sd-792, 8'sd65}},
{{13'sd2615, 12'sd1227, 13'sd2391}, {11'sd-818, 13'sd-2436, 11'sd-541}, {12'sd-1529, 11'sd-727, 12'sd-1904}}},
{
{{10'sd-264, 13'sd2805, 13'sd2401}, {12'sd-1238, 11'sd862, 13'sd-2244}, {12'sd-1654, 13'sd2111, 13'sd-3165}},
{{12'sd-1379, 10'sd-322, 13'sd2130}, {13'sd-2631, 6'sd-18, 12'sd-1150}, {8'sd-117, 13'sd-2991, 9'sd-178}},
{{12'sd1942, 9'sd251, 9'sd177}, {12'sd-1702, 12'sd1807, 13'sd2680}, {13'sd2089, 12'sd2025, 12'sd-1343}},
{{12'sd-1390, 13'sd2399, 11'sd995}, {9'sd128, 13'sd2535, 12'sd-1323}, {12'sd-1486, 13'sd-2335, 12'sd-1070}},
{{11'sd752, 11'sd-630, 7'sd56}, {12'sd-1143, 9'sd149, 13'sd-2606}, {11'sd-934, 10'sd392, 13'sd2176}},
{{5'sd12, 12'sd-1576, 12'sd-1539}, {13'sd2259, 11'sd801, 11'sd808}, {8'sd100, 12'sd-1123, 12'sd-1426}},
{{13'sd2906, 11'sd513, 12'sd2020}, {12'sd-1240, 12'sd-1213, 13'sd-2376}, {12'sd-1321, 6'sd-17, 13'sd-2075}},
{{12'sd1085, 10'sd-431, 13'sd2780}, {12'sd1927, 12'sd1096, 11'sd-602}, {13'sd-2493, 11'sd698, 12'sd-1295}},
{{12'sd1657, 12'sd-1433, 11'sd-723}, {12'sd1087, 12'sd1742, 12'sd1036}, {12'sd-1317, 6'sd-24, 13'sd2558}},
{{12'sd1210, 12'sd1320, 11'sd-617}, {13'sd-3144, 12'sd1470, 11'sd-755}, {13'sd-2422, 11'sd-630, 12'sd1285}},
{{14'sd4851, 7'sd49, 13'sd-3760}, {13'sd2272, 12'sd-2021, 8'sd-102}, {13'sd2048, 12'sd1245, 12'sd1164}},
{{12'sd-1617, 10'sd443, 12'sd1683}, {12'sd-1362, 12'sd1704, 11'sd-869}, {13'sd-2416, 13'sd-2541, 12'sd-1347}},
{{12'sd-1296, 11'sd637, 11'sd658}, {12'sd1830, 12'sd1958, 13'sd3441}, {12'sd-1140, 11'sd-517, 12'sd1453}},
{{12'sd-1683, 9'sd242, 9'sd-220}, {12'sd-1848, 12'sd1187, 11'sd-756}, {12'sd1043, 11'sd612, 13'sd2452}},
{{13'sd-2376, 12'sd-1806, 12'sd-1933}, {4'sd-5, 11'sd913, 12'sd-1371}, {12'sd-1916, 13'sd2335, 12'sd-1114}},
{{13'sd2365, 12'sd-1709, 13'sd3098}, {13'sd-2306, 13'sd2283, 12'sd-1115}, {12'sd1451, 12'sd1316, 10'sd-357}},
{{13'sd-2861, 11'sd-622, 12'sd-1081}, {11'sd973, 12'sd1796, 12'sd1960}, {12'sd1927, 13'sd2544, 11'sd-904}},
{{13'sd-3377, 11'sd646, 13'sd2049}, {12'sd-1393, 13'sd-2098, 12'sd1435}, {12'sd-2045, 12'sd1497, 11'sd655}},
{{13'sd2284, 13'sd2194, 11'sd934}, {13'sd2220, 13'sd-2077, 13'sd2262}, {12'sd1270, 11'sd-562, 10'sd405}},
{{13'sd2289, 11'sd965, 13'sd2262}, {10'sd445, 6'sd-18, 12'sd-1581}, {13'sd3045, 10'sd-328, 13'sd-2344}},
{{13'sd-2691, 13'sd-2630, 13'sd-2674}, {12'sd-2022, 8'sd-114, 12'sd-1205}, {11'sd-741, 13'sd-2411, 13'sd2371}},
{{13'sd-3203, 11'sd-959, 13'sd-2126}, {13'sd-2200, 12'sd1264, 10'sd-440}, {12'sd1661, 11'sd995, 12'sd1558}},
{{8'sd117, 13'sd-2775, 12'sd-1385}, {12'sd-1875, 13'sd-2777, 13'sd-2968}, {12'sd-1601, 12'sd-1409, 10'sd345}},
{{12'sd-1779, 11'sd897, 12'sd-1562}, {10'sd297, 12'sd1765, 9'sd229}, {12'sd-1947, 12'sd-1809, 12'sd-1524}},
{{12'sd-1480, 13'sd-3357, 8'sd116}, {8'sd93, 12'sd1723, 13'sd2256}, {13'sd-3067, 12'sd-1213, 13'sd2421}},
{{12'sd1893, 12'sd1030, 12'sd1856}, {12'sd1437, 13'sd2055, 12'sd-1056}, {12'sd-1277, 13'sd-2482, 8'sd-79}},
{{11'sd-889, 9'sd-221, 13'sd-2615}, {12'sd1081, 12'sd-1666, 11'sd856}, {8'sd112, 13'sd-2416, 12'sd1545}},
{{12'sd1271, 12'sd-1594, 12'sd1740}, {13'sd2164, 12'sd-1046, 12'sd1901}, {12'sd1878, 11'sd981, 8'sd103}},
{{8'sd80, 11'sd-878, 12'sd1036}, {12'sd1459, 13'sd2352, 11'sd-978}, {12'sd1428, 13'sd2328, 12'sd-1968}},
{{10'sd-324, 13'sd-2408, 11'sd-823}, {10'sd-508, 13'sd3120, 12'sd1471}, {13'sd2250, 11'sd-944, 13'sd2483}},
{{12'sd1469, 12'sd1461, 11'sd713}, {12'sd-1864, 12'sd1367, 11'sd-859}, {13'sd2489, 11'sd-972, 13'sd-2634}},
{{13'sd2908, 12'sd-1581, 7'sd-35}, {13'sd2366, 12'sd2017, 12'sd1037}, {13'sd-2049, 10'sd288, 13'sd-2644}},
{{13'sd-2332, 12'sd-2019, 13'sd2815}, {12'sd-1777, 8'sd126, 12'sd1282}, {13'sd-2519, 13'sd-2146, 12'sd1218}},
{{2'sd1, 12'sd-1596, 12'sd-1050}, {13'sd2454, 13'sd2134, 12'sd-1983}, {11'sd837, 11'sd606, 12'sd-1674}},
{{11'sd1022, 10'sd479, 10'sd286}, {13'sd2365, 12'sd1860, 11'sd-564}, {12'sd1131, 13'sd-2584, 10'sd317}},
{{12'sd-1952, 10'sd505, 13'sd-2774}, {10'sd272, 12'sd1658, 9'sd-132}, {13'sd-2481, 13'sd2691, 11'sd724}},
{{11'sd-608, 10'sd384, 13'sd2298}, {13'sd-2447, 11'sd-987, 12'sd1185}, {13'sd-2181, 12'sd-1307, 11'sd-1003}},
{{12'sd-1333, 13'sd2687, 12'sd-1874}, {12'sd-1829, 12'sd-1743, 12'sd1655}, {12'sd-1173, 11'sd953, 11'sd-846}},
{{11'sd-770, 12'sd1863, 13'sd2236}, {13'sd-2915, 12'sd-1612, 11'sd792}, {9'sd169, 11'sd587, 11'sd551}},
{{11'sd-780, 12'sd1336, 11'sd-581}, {11'sd-744, 13'sd2101, 12'sd-1987}, {13'sd-2568, 13'sd-2173, 10'sd-320}},
{{11'sd-900, 13'sd2334, 12'sd2021}, {12'sd1066, 12'sd1217, 12'sd1071}, {13'sd-2411, 10'sd446, 8'sd96}},
{{12'sd-1119, 11'sd728, 12'sd1656}, {13'sd2063, 12'sd1616, 9'sd159}, {13'sd-2435, 12'sd1633, 12'sd1980}},
{{12'sd1647, 11'sd720, 10'sd494}, {12'sd-1723, 12'sd-1080, 13'sd-2476}, {12'sd1807, 12'sd-1418, 13'sd2153}},
{{12'sd-1834, 13'sd2253, 11'sd847}, {12'sd1047, 12'sd-1405, 11'sd519}, {12'sd1206, 12'sd-1779, 13'sd2289}},
{{13'sd-2485, 12'sd1544, 12'sd1037}, {11'sd-749, 9'sd169, 11'sd687}, {13'sd-2247, 11'sd812, 12'sd1882}},
{{13'sd-2921, 13'sd-2819, 12'sd1693}, {12'sd-1892, 11'sd945, 13'sd2308}, {12'sd1904, 9'sd-198, 8'sd72}},
{{12'sd-1548, 12'sd1393, 12'sd1443}, {11'sd-767, 12'sd-1931, 11'sd-572}, {6'sd22, 9'sd142, 12'sd-1978}},
{{13'sd2412, 13'sd2270, 11'sd872}, {12'sd-1238, 12'sd-1070, 10'sd383}, {12'sd1767, 11'sd-646, 11'sd-762}},
{{11'sd-662, 10'sd-340, 7'sd-63}, {10'sd-448, 12'sd-1644, 10'sd-463}, {10'sd-436, 8'sd-88, 11'sd669}},
{{12'sd-1308, 10'sd-430, 11'sd-682}, {13'sd2264, 10'sd-484, 13'sd2370}, {11'sd702, 13'sd2434, 12'sd-1587}},
{{13'sd2203, 13'sd2401, 11'sd872}, {9'sd241, 11'sd-860, 12'sd1215}, {12'sd-1564, 10'sd-339, 12'sd-1962}},
{{3'sd-3, 12'sd-1036, 11'sd895}, {12'sd1747, 12'sd1979, 12'sd1203}, {13'sd2323, 12'sd-1232, 13'sd-2138}},
{{12'sd-1820, 13'sd-2757, 12'sd1367}, {13'sd-2403, 9'sd240, 13'sd-3551}, {13'sd-2313, 10'sd-468, 11'sd-741}},
{{13'sd-2391, 13'sd2147, 13'sd2779}, {12'sd-1685, 10'sd-285, 12'sd1172}, {11'sd-1013, 12'sd1236, 9'sd163}},
{{12'sd1768, 13'sd2342, 11'sd-716}, {12'sd-1964, 12'sd-1405, 11'sd575}, {10'sd-465, 13'sd-3006, 12'sd-1683}},
{{10'sd-355, 13'sd-2595, 9'sd212}, {10'sd-334, 10'sd439, 12'sd1637}, {12'sd-1867, 9'sd215, 13'sd-2378}},
{{13'sd2676, 13'sd2052, 12'sd1861}, {11'sd-993, 12'sd1284, 10'sd-379}, {12'sd-1325, 13'sd-2480, 11'sd-856}},
{{13'sd2072, 13'sd2547, 11'sd-980}, {11'sd-964, 12'sd-1099, 11'sd-978}, {12'sd-1917, 13'sd2297, 10'sd350}},
{{12'sd1396, 11'sd1009, 11'sd951}, {12'sd1670, 13'sd-2889, 12'sd1031}, {11'sd-853, 12'sd1844, 11'sd896}},
{{13'sd-2722, 11'sd-884, 13'sd-2250}, {12'sd-1056, 11'sd702, 12'sd1093}, {13'sd2258, 12'sd-1185, 7'sd60}},
{{13'sd-2423, 10'sd259, 13'sd-2342}, {11'sd763, 13'sd2677, 12'sd1614}, {10'sd-478, 12'sd-1972, 9'sd253}},
{{12'sd-1243, 13'sd2240, 12'sd-1626}, {10'sd340, 12'sd1375, 12'sd1990}, {12'sd-1038, 12'sd-1406, 6'sd29}},
{{12'sd-1946, 11'sd648, 10'sd327}, {12'sd1496, 12'sd1313, 12'sd-1567}, {8'sd102, 12'sd1996, 12'sd1304}},
{{13'sd-3019, 8'sd88, 12'sd1423}, {12'sd1931, 12'sd-1711, 13'sd-2844}, {12'sd-1820, 12'sd-1902, 11'sd-709}}},
{
{{13'sd-2889, 12'sd-1809, 12'sd1029}, {10'sd303, 11'sd607, 9'sd-144}, {11'sd546, 12'sd1347, 13'sd-2301}},
{{9'sd-138, 12'sd1477, 12'sd1623}, {8'sd-64, 11'sd-594, 11'sd-704}, {13'sd-3138, 12'sd1073, 12'sd-1400}},
{{14'sd4805, 13'sd-2923, 11'sd556}, {12'sd1698, 13'sd-3863, 12'sd1699}, {13'sd2694, 9'sd-248, 10'sd494}},
{{11'sd1003, 13'sd2070, 12'sd1299}, {12'sd1809, 11'sd695, 12'sd1921}, {12'sd-1625, 13'sd2174, 12'sd1542}},
{{12'sd-1110, 13'sd2441, 12'sd1668}, {10'sd334, 12'sd1640, 9'sd229}, {13'sd-2807, 12'sd1836, 11'sd553}},
{{10'sd-493, 5'sd-13, 13'sd-3097}, {12'sd1137, 12'sd-1555, 12'sd1903}, {12'sd-1448, 10'sd468, 13'sd-2269}},
{{12'sd1637, 10'sd485, 13'sd-2576}, {11'sd586, 12'sd-1921, 12'sd1408}, {11'sd-553, 11'sd538, 11'sd626}},
{{13'sd-2486, 13'sd-2262, 12'sd-1718}, {12'sd1467, 11'sd-725, 11'sd777}, {13'sd4000, 9'sd-140, 12'sd1410}},
{{12'sd-1239, 12'sd-1971, 12'sd2038}, {11'sd-890, 12'sd1363, 12'sd-1071}, {12'sd-1444, 13'sd2307, 11'sd-808}},
{{12'sd1056, 11'sd668, 12'sd-1981}, {13'sd-2060, 10'sd469, 12'sd1982}, {11'sd655, 13'sd-2198, 11'sd-537}},
{{12'sd-1132, 13'sd-2602, 14'sd-4785}, {12'sd-1078, 12'sd1145, 12'sd-1897}, {12'sd1137, 13'sd2403, 13'sd2280}},
{{12'sd-1342, 13'sd2720, 8'sd-68}, {12'sd1956, 12'sd2000, 12'sd1136}, {13'sd2830, 13'sd-2101, 13'sd2998}},
{{12'sd1755, 13'sd-2795, 12'sd1244}, {12'sd-1627, 13'sd-3127, 10'sd-450}, {12'sd-1183, 13'sd2104, 11'sd540}},
{{11'sd-805, 13'sd2900, 12'sd-1956}, {11'sd667, 13'sd-2335, 11'sd852}, {10'sd353, 13'sd2137, 13'sd2300}},
{{12'sd1648, 12'sd1369, 7'sd55}, {11'sd-574, 12'sd-1829, 10'sd-463}, {13'sd-2210, 12'sd1536, 12'sd1366}},
{{12'sd-1493, 11'sd891, 12'sd-1583}, {8'sd-124, 12'sd-1285, 13'sd2176}, {13'sd2420, 12'sd-1255, 12'sd-1715}},
{{13'sd-3374, 13'sd-2504, 11'sd978}, {11'sd-776, 12'sd-1178, 13'sd2996}, {12'sd1461, 13'sd-3056, 12'sd1813}},
{{14'sd4866, 13'sd2294, 13'sd2563}, {12'sd-1401, 13'sd2098, 13'sd-2108}, {9'sd-145, 11'sd-1006, 13'sd-2447}},
{{13'sd2419, 10'sd318, 13'sd2302}, {12'sd-1933, 11'sd977, 12'sd-1866}, {13'sd2644, 13'sd-2273, 11'sd-816}},
{{12'sd1156, 11'sd788, 11'sd-529}, {12'sd1543, 13'sd3073, 8'sd-79}, {12'sd-1930, 13'sd2753, 12'sd-1120}},
{{12'sd1044, 12'sd1686, 13'sd-3118}, {13'sd2695, 12'sd1223, 13'sd-2149}, {12'sd1459, 12'sd-1648, 10'sd-421}},
{{13'sd3068, 9'sd-238, 12'sd-1665}, {11'sd986, 13'sd-3736, 12'sd-1650}, {9'sd203, 11'sd-1004, 13'sd-3062}},
{{13'sd2752, 13'sd-2240, 12'sd1333}, {12'sd1246, 11'sd-654, 13'sd-2205}, {12'sd-1169, 13'sd2128, 11'sd640}},
{{11'sd-600, 13'sd2818, 12'sd1206}, {13'sd2609, 12'sd-1120, 13'sd-3166}, {11'sd-759, 13'sd2164, 11'sd-738}},
{{13'sd3093, 12'sd-1836, 12'sd1768}, {11'sd-685, 12'sd-1268, 11'sd649}, {12'sd-1374, 13'sd-3832, 13'sd2192}},
{{12'sd2003, 13'sd2664, 11'sd813}, {12'sd1047, 12'sd1655, 12'sd-1206}, {12'sd-1872, 12'sd-1684, 11'sd785}},
{{10'sd314, 13'sd2134, 13'sd3282}, {12'sd1513, 11'sd-631, 12'sd-1481}, {11'sd836, 12'sd-1488, 13'sd2335}},
{{12'sd-1798, 9'sd128, 11'sd990}, {12'sd1056, 13'sd-2055, 12'sd1092}, {13'sd-2463, 11'sd1009, 10'sd-458}},
{{12'sd-1086, 11'sd-706, 12'sd1855}, {12'sd-1517, 13'sd-2376, 10'sd338}, {12'sd-1452, 13'sd-2378, 8'sd115}},
{{13'sd-3438, 14'sd-4643, 13'sd2872}, {10'sd-482, 13'sd-2456, 12'sd-1304}, {13'sd-2717, 10'sd-442, 9'sd148}},
{{11'sd-796, 12'sd-1194, 13'sd-2294}, {12'sd1634, 11'sd567, 12'sd1028}, {13'sd-2717, 12'sd-1099, 11'sd556}},
{{12'sd-1688, 12'sd-1634, 12'sd1324}, {13'sd2407, 13'sd2885, 12'sd1524}, {11'sd-721, 11'sd1007, 13'sd-3074}},
{{11'sd1007, 12'sd-1112, 13'sd-2114}, {11'sd-928, 8'sd87, 12'sd-1761}, {12'sd1817, 10'sd427, 12'sd1148}},
{{12'sd-1275, 13'sd-2500, 13'sd-2365}, {10'sd-358, 12'sd-1144, 10'sd-386}, {13'sd2229, 8'sd113, 12'sd1638}},
{{13'sd-2459, 10'sd403, 12'sd-1988}, {12'sd-1055, 11'sd-860, 13'sd2120}, {11'sd953, 8'sd-115, 13'sd-2523}},
{{11'sd-956, 12'sd1170, 13'sd2647}, {11'sd-915, 12'sd-1555, 13'sd2500}, {12'sd-1601, 12'sd-1176, 13'sd2858}},
{{8'sd97, 13'sd2857, 11'sd-1003}, {13'sd2550, 12'sd-1791, 8'sd-109}, {11'sd520, 12'sd1637, 13'sd2196}},
{{14'sd-4707, 13'sd-2422, 11'sd727}, {13'sd-2714, 10'sd-378, 9'sd-249}, {12'sd-1728, 9'sd-135, 13'sd3088}},
{{10'sd-315, 12'sd-1777, 11'sd-856}, {12'sd-2020, 9'sd-134, 9'sd143}, {12'sd-1752, 13'sd2972, 11'sd-753}},
{{11'sd644, 13'sd2601, 12'sd-1744}, {9'sd214, 13'sd2308, 12'sd-1775}, {11'sd598, 11'sd-686, 12'sd-1856}},
{{12'sd1161, 12'sd1199, 13'sd-3592}, {12'sd1895, 11'sd702, 12'sd1622}, {13'sd-2522, 13'sd-2729, 12'sd-1912}},
{{12'sd1980, 13'sd-2135, 12'sd1622}, {12'sd-1293, 7'sd-62, 12'sd-1170}, {12'sd-1515, 10'sd-332, 12'sd-1869}},
{{11'sd-701, 13'sd3534, 11'sd-1007}, {9'sd173, 12'sd1256, 12'sd1217}, {8'sd103, 12'sd1037, 9'sd252}},
{{11'sd-772, 11'sd534, 11'sd-561}, {13'sd-2464, 10'sd330, 11'sd982}, {11'sd-530, 12'sd1309, 13'sd2393}},
{{12'sd1962, 10'sd-437, 9'sd-155}, {9'sd-255, 13'sd-2484, 11'sd-748}, {11'sd-526, 13'sd-2885, 12'sd1852}},
{{13'sd2993, 13'sd2166, 13'sd-2523}, {12'sd1430, 13'sd2590, 11'sd759}, {9'sd180, 13'sd-2197, 12'sd1713}},
{{12'sd1557, 11'sd-617, 12'sd1862}, {12'sd-1764, 12'sd-1378, 13'sd3155}, {12'sd1735, 13'sd2172, 13'sd-2476}},
{{12'sd1939, 12'sd1932, 13'sd-3296}, {12'sd-1131, 12'sd-1615, 11'sd884}, {12'sd-1714, 12'sd1847, 12'sd1214}},
{{12'sd-1131, 13'sd2490, 11'sd-819}, {7'sd-35, 8'sd120, 13'sd2217}, {11'sd798, 12'sd-1163, 9'sd137}},
{{12'sd-1596, 10'sd294, 11'sd972}, {9'sd177, 12'sd-1510, 11'sd790}, {12'sd1253, 12'sd-1982, 12'sd1219}},
{{13'sd2358, 12'sd-1453, 10'sd-510}, {13'sd-2593, 11'sd773, 11'sd-864}, {9'sd-135, 12'sd-1959, 13'sd3034}},
{{13'sd2386, 12'sd-1984, 12'sd-1404}, {13'sd-2251, 13'sd-2387, 11'sd762}, {13'sd2560, 7'sd52, 11'sd-837}},
{{12'sd1155, 12'sd-1225, 13'sd-2685}, {9'sd225, 12'sd1970, 11'sd-579}, {11'sd-680, 9'sd-160, 11'sd-714}},
{{12'sd1849, 13'sd2740, 11'sd-619}, {11'sd-673, 12'sd1132, 12'sd1610}, {12'sd1436, 10'sd-425, 13'sd2163}},
{{11'sd-810, 13'sd2475, 12'sd1318}, {13'sd2115, 12'sd1116, 9'sd237}, {12'sd1348, 12'sd-1863, 11'sd556}},
{{12'sd-1749, 13'sd2105, 10'sd-490}, {12'sd1415, 10'sd-496, 11'sd797}, {13'sd2120, 8'sd81, 12'sd-1849}},
{{13'sd2098, 11'sd711, 9'sd154}, {12'sd1463, 13'sd-2448, 13'sd-2547}, {13'sd2632, 12'sd-1774, 12'sd1158}},
{{13'sd-2181, 11'sd-513, 11'sd517}, {10'sd-406, 12'sd1789, 11'sd-863}, {13'sd2809, 12'sd1131, 11'sd-795}},
{{13'sd2709, 12'sd1154, 12'sd1566}, {11'sd-897, 13'sd2154, 12'sd-1891}, {12'sd-1436, 7'sd-37, 12'sd-1304}},
{{13'sd-2492, 11'sd-625, 11'sd604}, {13'sd-2198, 11'sd-970, 9'sd233}, {10'sd406, 12'sd1750, 11'sd853}},
{{13'sd-2203, 12'sd-1090, 13'sd3253}, {12'sd1949, 8'sd-80, 13'sd2862}, {12'sd1774, 13'sd-3086, 10'sd382}},
{{8'sd-77, 13'sd2064, 9'sd224}, {8'sd94, 10'sd-476, 12'sd-1192}, {13'sd2495, 9'sd205, 10'sd377}},
{{13'sd-2337, 12'sd1667, 11'sd-618}, {12'sd-1750, 12'sd-1408, 11'sd-543}, {12'sd1311, 11'sd-579, 12'sd-1668}},
{{9'sd-143, 9'sd-135, 13'sd2599}, {13'sd-2672, 13'sd-2841, 10'sd-351}, {12'sd-1647, 13'sd2322, 9'sd201}}},
{
{{13'sd2520, 11'sd639, 13'sd2225}, {13'sd-2543, 13'sd-2246, 13'sd-3172}, {13'sd-2660, 13'sd-3345, 13'sd-3555}},
{{13'sd-3089, 11'sd689, 10'sd306}, {11'sd884, 12'sd-1459, 13'sd2150}, {13'sd-2669, 8'sd-75, 11'sd-1022}},
{{12'sd1842, 12'sd1197, 12'sd1649}, {12'sd-1891, 13'sd-2638, 10'sd-329}, {12'sd-1878, 12'sd1383, 12'sd1737}},
{{13'sd-2357, 12'sd-1107, 12'sd-1827}, {13'sd2455, 8'sd93, 12'sd-1200}, {12'sd-1997, 12'sd1557, 13'sd-2246}},
{{8'sd-121, 13'sd-2253, 12'sd-1065}, {12'sd-1941, 13'sd-2747, 12'sd1932}, {12'sd-1504, 11'sd-936, 12'sd1129}},
{{13'sd2446, 12'sd-1919, 13'sd2497}, {10'sd-417, 11'sd732, 11'sd908}, {12'sd-1585, 13'sd-2539, 12'sd-1114}},
{{10'sd286, 11'sd-653, 12'sd1270}, {12'sd-1904, 12'sd1834, 12'sd1085}, {13'sd2193, 13'sd2057, 12'sd-1060}},
{{13'sd2207, 12'sd1288, 12'sd1934}, {12'sd1089, 9'sd135, 12'sd-1460}, {12'sd1273, 12'sd-1396, 12'sd-1969}},
{{12'sd1862, 11'sd777, 11'sd-615}, {13'sd-2143, 10'sd304, 12'sd1605}, {13'sd2881, 9'sd-155, 13'sd-2237}},
{{5'sd-11, 13'sd2276, 12'sd-1282}, {11'sd940, 12'sd1936, 13'sd2126}, {12'sd-1561, 13'sd-2288, 11'sd-746}},
{{12'sd-1062, 11'sd-642, 11'sd902}, {13'sd-2470, 12'sd1976, 11'sd-871}, {13'sd2619, 14'sd4185, 13'sd3771}},
{{12'sd1092, 9'sd135, 11'sd-886}, {11'sd790, 13'sd-2864, 8'sd-94}, {13'sd-2103, 13'sd2689, 12'sd1137}},
{{9'sd241, 11'sd-788, 13'sd2870}, {13'sd-3041, 10'sd310, 11'sd939}, {12'sd1801, 9'sd-184, 11'sd984}},
{{12'sd1108, 9'sd244, 12'sd1932}, {9'sd128, 13'sd-2253, 7'sd-33}, {12'sd-1346, 13'sd-2108, 12'sd1535}},
{{13'sd-2136, 12'sd1578, 12'sd1437}, {7'sd44, 12'sd1748, 13'sd-2490}, {13'sd2201, 11'sd-848, 11'sd-980}},
{{13'sd2098, 11'sd1006, 11'sd874}, {12'sd1384, 13'sd-2415, 12'sd-1501}, {10'sd-487, 10'sd-261, 10'sd283}},
{{12'sd1658, 13'sd2183, 11'sd-518}, {12'sd1082, 12'sd-1442, 12'sd1799}, {13'sd-2569, 8'sd-114, 12'sd-2035}},
{{13'sd4074, 12'sd1443, 13'sd2228}, {13'sd2719, 13'sd2530, 13'sd2984}, {13'sd2194, 13'sd2070, 13'sd2269}},
{{12'sd-1744, 11'sd965, 13'sd3101}, {10'sd325, 11'sd599, 11'sd1017}, {12'sd1134, 13'sd-2060, 10'sd318}},
{{13'sd3084, 13'sd3146, 11'sd-807}, {11'sd-1018, 12'sd-1506, 13'sd2655}, {8'sd105, 12'sd1475, 12'sd-1740}},
{{13'sd2446, 13'sd2782, 12'sd1637}, {13'sd-2259, 11'sd-915, 10'sd470}, {12'sd1453, 11'sd-974, 9'sd-246}},
{{12'sd-1707, 13'sd-2787, 12'sd-1413}, {13'sd-2908, 12'sd-1691, 13'sd-3759}, {12'sd-1523, 12'sd-1878, 11'sd-815}},
{{9'sd-172, 9'sd135, 13'sd-3235}, {11'sd763, 12'sd-1932, 12'sd1377}, {10'sd282, 13'sd2247, 11'sd936}},
{{12'sd1906, 13'sd2187, 11'sd869}, {12'sd-1443, 13'sd-2706, 11'sd599}, {12'sd-1284, 11'sd745, 13'sd2710}},
{{13'sd-2608, 9'sd-213, 12'sd-1899}, {3'sd-2, 12'sd-1970, 12'sd-1568}, {11'sd-982, 13'sd-3301, 11'sd-803}},
{{11'sd913, 13'sd2816, 12'sd-1241}, {12'sd-1465, 11'sd-586, 13'sd2424}, {13'sd-2232, 11'sd-927, 12'sd-1206}},
{{13'sd2253, 13'sd2320, 11'sd733}, {9'sd-192, 12'sd1731, 12'sd1593}, {6'sd-30, 12'sd-1746, 11'sd929}},
{{13'sd3058, 13'sd2287, 11'sd738}, {13'sd3226, 11'sd-930, 10'sd-369}, {6'sd-30, 12'sd-1515, 11'sd-564}},
{{13'sd2368, 13'sd-2227, 11'sd-587}, {12'sd-1488, 10'sd469, 12'sd1908}, {9'sd176, 13'sd2605, 12'sd-1067}},
{{10'sd457, 12'sd-1919, 11'sd684}, {11'sd829, 12'sd-1746, 6'sd27}, {12'sd-1119, 13'sd-2583, 11'sd691}},
{{12'sd1989, 13'sd-2762, 12'sd-1475}, {12'sd-1549, 11'sd-668, 12'sd1362}, {11'sd571, 9'sd251, 6'sd28}},
{{12'sd-1698, 12'sd-1822, 12'sd-1531}, {12'sd-1874, 12'sd1383, 11'sd949}, {11'sd519, 12'sd-1892, 13'sd-2424}},
{{11'sd-863, 12'sd1288, 12'sd1197}, {10'sd436, 10'sd479, 12'sd-1436}, {12'sd1039, 10'sd-428, 11'sd-765}},
{{12'sd1731, 11'sd586, 10'sd508}, {12'sd-1412, 11'sd739, 13'sd2096}, {12'sd1982, 13'sd2656, 12'sd-1201}},
{{10'sd-497, 12'sd-1797, 12'sd-1343}, {13'sd2370, 13'sd2244, 9'sd-248}, {12'sd1959, 10'sd434, 12'sd1565}},
{{11'sd-890, 11'sd-785, 12'sd1284}, {12'sd-1599, 13'sd-2302, 13'sd2148}, {12'sd1150, 10'sd-431, 13'sd-2154}},
{{12'sd1817, 13'sd2615, 12'sd1394}, {12'sd1631, 13'sd-2753, 10'sd340}, {12'sd1946, 12'sd-1738, 10'sd349}},
{{11'sd-629, 13'sd-3278, 13'sd2645}, {10'sd-305, 13'sd-3109, 12'sd1849}, {8'sd-70, 13'sd-2058, 12'sd-1256}},
{{12'sd1860, 11'sd-716, 12'sd-1611}, {10'sd-466, 11'sd-900, 11'sd-839}, {11'sd-705, 12'sd1731, 11'sd-905}},
{{12'sd-1387, 10'sd-490, 10'sd-352}, {12'sd-1234, 13'sd2545, 12'sd-1939}, {11'sd-619, 10'sd-302, 12'sd-1354}},
{{10'sd-468, 12'sd1255, 9'sd154}, {11'sd558, 6'sd-19, 12'sd1155}, {13'sd-3001, 11'sd987, 12'sd-1456}},
{{13'sd2684, 12'sd1749, 10'sd494}, {13'sd-2308, 12'sd1536, 12'sd2009}, {13'sd2127, 12'sd-1309, 11'sd-550}},
{{12'sd-1115, 13'sd-2386, 9'sd-190}, {11'sd-791, 11'sd909, 11'sd-919}, {12'sd-1078, 11'sd748, 12'sd-1948}},
{{12'sd1129, 7'sd46, 11'sd848}, {13'sd2179, 11'sd-828, 11'sd-766}, {8'sd-94, 9'sd-154, 11'sd-651}},
{{11'sd-1005, 12'sd-1286, 12'sd1083}, {10'sd-397, 12'sd1093, 12'sd-1928}, {11'sd963, 11'sd830, 12'sd-1946}},
{{12'sd1044, 11'sd-648, 5'sd11}, {13'sd-2085, 10'sd-494, 11'sd933}, {12'sd-1699, 12'sd2001, 12'sd-1788}},
{{10'sd473, 12'sd1161, 6'sd-30}, {13'sd2259, 7'sd32, 9'sd133}, {12'sd-1066, 12'sd1861, 12'sd-1159}},
{{10'sd-485, 12'sd2006, 12'sd-1512}, {6'sd30, 12'sd1933, 8'sd111}, {13'sd-3067, 12'sd1221, 12'sd1764}},
{{13'sd2297, 11'sd837, 13'sd-2355}, {13'sd2412, 13'sd-2160, 11'sd-770}, {10'sd-264, 12'sd-1398, 12'sd-1562}},
{{12'sd1221, 12'sd-1596, 11'sd-846}, {11'sd-1005, 12'sd-1810, 10'sd317}, {12'sd1738, 12'sd1721, 12'sd-1426}},
{{11'sd-888, 12'sd1414, 13'sd2242}, {10'sd375, 13'sd-2220, 9'sd-164}, {12'sd1465, 13'sd2534, 12'sd1426}},
{{13'sd3285, 11'sd-1002, 12'sd-1399}, {13'sd2937, 12'sd-2042, 12'sd-1699}, {11'sd-647, 13'sd2549, 13'sd-2257}},
{{12'sd1158, 13'sd-2651, 11'sd851}, {12'sd-1733, 12'sd-1274, 9'sd224}, {12'sd-1585, 9'sd154, 10'sd-449}},
{{12'sd1623, 10'sd330, 13'sd-3051}, {12'sd1834, 13'sd-2788, 13'sd2422}, {13'sd-2332, 10'sd263, 13'sd2293}},
{{13'sd-2960, 12'sd1261, 11'sd696}, {10'sd370, 13'sd-2183, 11'sd905}, {12'sd-1027, 12'sd1802, 13'sd2273}},
{{11'sd613, 10'sd326, 13'sd2740}, {12'sd-1767, 8'sd102, 10'sd451}, {13'sd2405, 13'sd2397, 12'sd1658}},
{{12'sd1335, 12'sd-1695, 11'sd792}, {13'sd-2707, 12'sd-1065, 9'sd158}, {12'sd-1631, 13'sd3002, 9'sd202}},
{{11'sd-525, 12'sd-1882, 13'sd2286}, {13'sd3102, 12'sd-1196, 5'sd11}, {11'sd-771, 13'sd2578, 12'sd1581}},
{{12'sd-1803, 12'sd-1746, 13'sd-3298}, {12'sd1211, 12'sd-1680, 13'sd2283}, {13'sd2863, 13'sd-2585, 9'sd131}},
{{12'sd1480, 11'sd798, 13'sd2443}, {13'sd-2356, 12'sd1997, 12'sd1823}, {11'sd-970, 12'sd1559, 11'sd-942}},
{{11'sd624, 12'sd-1634, 11'sd-705}, {13'sd2255, 13'sd-2089, 12'sd1535}, {9'sd211, 12'sd-1397, 12'sd-1632}},
{{11'sd-997, 13'sd2614, 12'sd1794}, {11'sd-535, 12'sd1696, 10'sd-416}, {12'sd1457, 12'sd-1635, 11'sd689}},
{{13'sd-2489, 13'sd2411, 9'sd-184}, {11'sd-726, 11'sd675, 8'sd-93}, {12'sd-1837, 12'sd-1855, 11'sd-837}},
{{10'sd369, 12'sd1892, 13'sd2565}, {12'sd-1447, 12'sd-1370, 11'sd-779}, {13'sd-2910, 12'sd-1374, 12'sd1830}}},
{
{{11'sd994, 11'sd529, 12'sd1061}, {11'sd-523, 12'sd-1870, 12'sd1294}, {11'sd-525, 10'sd-499, 10'sd-492}},
{{12'sd1661, 9'sd-177, 12'sd1986}, {12'sd-1843, 13'sd2756, 12'sd1367}, {13'sd-3830, 13'sd3007, 12'sd1358}},
{{13'sd-3260, 11'sd-552, 12'sd1296}, {12'sd-1873, 13'sd2914, 12'sd1071}, {13'sd-3624, 13'sd2479, 13'sd2322}},
{{9'sd-190, 12'sd-1177, 11'sd-630}, {13'sd3005, 9'sd213, 12'sd1276}, {13'sd2954, 12'sd-1321, 11'sd-885}},
{{13'sd3794, 13'sd2890, 13'sd-2061}, {13'sd2290, 13'sd2410, 12'sd1943}, {12'sd1220, 10'sd-289, 11'sd730}},
{{13'sd-2129, 13'sd-2886, 11'sd984}, {12'sd-1727, 12'sd-1305, 12'sd1426}, {12'sd1475, 13'sd-2691, 12'sd1064}},
{{8'sd116, 10'sd377, 12'sd-1804}, {13'sd-2814, 13'sd-3387, 13'sd-3953}, {13'sd-2875, 10'sd279, 13'sd-3337}},
{{13'sd3042, 9'sd248, 13'sd3186}, {12'sd1411, 11'sd-855, 13'sd-2166}, {10'sd-332, 12'sd1198, 10'sd389}},
{{13'sd-2095, 11'sd-611, 12'sd-1539}, {12'sd1498, 12'sd1361, 12'sd1812}, {10'sd439, 13'sd2314, 12'sd1465}},
{{12'sd1652, 6'sd30, 13'sd-2751}, {13'sd-3646, 8'sd86, 13'sd-2230}, {13'sd-3390, 12'sd-1840, 13'sd-2656}},
{{14'sd-4342, 12'sd-1489, 13'sd-3019}, {12'sd1786, 10'sd386, 12'sd1295}, {13'sd-3236, 8'sd109, 12'sd-1755}},
{{11'sd-926, 12'sd1541, 11'sd996}, {12'sd-1180, 11'sd-528, 12'sd-1294}, {12'sd1138, 13'sd2705, 13'sd2143}},
{{12'sd1717, 14'sd5174, 14'sd4247}, {11'sd-965, 12'sd1595, 12'sd-1707}, {10'sd-434, 9'sd227, 12'sd1671}},
{{12'sd1280, 13'sd-2366, 12'sd1451}, {12'sd-1790, 12'sd-1577, 9'sd-134}, {13'sd3293, 6'sd23, 10'sd393}},
{{13'sd2070, 12'sd-1697, 11'sd618}, {13'sd-2831, 11'sd-771, 9'sd245}, {13'sd-3512, 12'sd-1458, 11'sd-852}},
{{9'sd-144, 12'sd1043, 10'sd503}, {13'sd2935, 12'sd1835, 12'sd1883}, {12'sd-1152, 11'sd707, 13'sd-2683}},
{{13'sd-2204, 11'sd959, 12'sd-1465}, {11'sd-532, 13'sd3414, 13'sd3131}, {10'sd-349, 9'sd-218, 13'sd-2404}},
{{10'sd-313, 13'sd-2541, 12'sd1206}, {14'sd-4192, 9'sd-231, 11'sd-922}, {13'sd-2394, 14'sd-4743, 14'sd-5394}},
{{11'sd-881, 13'sd-2206, 10'sd-417}, {11'sd-688, 11'sd930, 12'sd1477}, {11'sd807, 11'sd-982, 12'sd-1648}},
{{13'sd2765, 13'sd2570, 9'sd-252}, {11'sd-762, 11'sd671, 12'sd1172}, {13'sd-2954, 12'sd-1579, 12'sd-1710}},
{{14'sd-4864, 12'sd-1707, 12'sd1046}, {10'sd324, 12'sd-1344, 13'sd2242}, {12'sd-1691, 12'sd1340, 12'sd1059}},
{{11'sd-628, 9'sd219, 12'sd1660}, {13'sd2254, 13'sd2857, 12'sd-1889}, {13'sd-3875, 11'sd560, 12'sd-1087}},
{{11'sd727, 9'sd-160, 12'sd-1377}, {11'sd782, 11'sd-870, 10'sd-427}, {10'sd-502, 12'sd1172, 10'sd387}},
{{11'sd-766, 11'sd-857, 12'sd-1470}, {11'sd666, 8'sd103, 11'sd-671}, {9'sd212, 9'sd205, 12'sd-1157}},
{{12'sd1208, 11'sd995, 13'sd2433}, {12'sd1333, 12'sd1595, 11'sd538}, {13'sd3974, 14'sd5440, 14'sd6003}},
{{9'sd200, 11'sd691, 12'sd-1751}, {13'sd2337, 12'sd1158, 12'sd-1685}, {12'sd-1675, 7'sd37, 7'sd-35}},
{{12'sd1524, 12'sd1451, 12'sd-1834}, {12'sd1117, 11'sd648, 11'sd727}, {13'sd2357, 10'sd483, 13'sd-2447}},
{{12'sd1770, 11'sd-750, 13'sd-2335}, {8'sd70, 11'sd781, 13'sd-3293}, {13'sd-2491, 12'sd-1607, 11'sd-682}},
{{9'sd-167, 12'sd-1725, 10'sd-449}, {12'sd1922, 10'sd-501, 11'sd-652}, {9'sd227, 12'sd-1960, 11'sd899}},
{{12'sd1328, 12'sd-1164, 10'sd-323}, {11'sd697, 8'sd-123, 13'sd-3168}, {13'sd-2459, 13'sd-2221, 12'sd1158}},
{{13'sd2844, 12'sd1570, 12'sd-1871}, {9'sd148, 13'sd2295, 13'sd3170}, {13'sd-2212, 12'sd1341, 11'sd1009}},
{{8'sd-68, 12'sd1928, 11'sd-575}, {11'sd612, 12'sd-1118, 12'sd-1826}, {3'sd2, 14'sd-4543, 11'sd836}},
{{13'sd-2645, 12'sd-1516, 13'sd2442}, {13'sd-2311, 12'sd1845, 10'sd-325}, {12'sd-1791, 13'sd-2390, 13'sd-2691}},
{{12'sd-1828, 13'sd2301, 12'sd1336}, {12'sd-1543, 12'sd1327, 12'sd1794}, {13'sd3009, 12'sd1868, 11'sd-672}},
{{12'sd1048, 12'sd1637, 10'sd-461}, {11'sd695, 12'sd1215, 13'sd2149}, {12'sd1207, 11'sd858, 12'sd-1979}},
{{13'sd2863, 12'sd-1443, 12'sd1964}, {12'sd-1708, 10'sd337, 10'sd-321}, {12'sd1549, 12'sd1251, 12'sd-1592}},
{{13'sd-2065, 13'sd-2068, 11'sd953}, {11'sd563, 13'sd2310, 12'sd1847}, {13'sd-3134, 11'sd-600, 13'sd2190}},
{{12'sd1062, 13'sd2827, 13'sd2590}, {14'sd4604, 13'sd-2318, 12'sd-1246}, {13'sd-3792, 13'sd-3485, 13'sd-2928}},
{{13'sd-2811, 11'sd-955, 14'sd6088}, {8'sd114, 10'sd258, 11'sd850}, {13'sd-2745, 11'sd-984, 13'sd2081}},
{{13'sd-2692, 13'sd3306, 13'sd3398}, {12'sd-1999, 13'sd-2103, 13'sd2872}, {13'sd-4054, 8'sd111, 13'sd-2429}},
{{11'sd692, 11'sd-900, 13'sd3498}, {7'sd-56, 12'sd1054, 13'sd3279}, {13'sd2092, 10'sd275, 12'sd-1492}},
{{13'sd2329, 12'sd-1822, 12'sd-1221}, {11'sd-849, 10'sd374, 13'sd-2680}, {10'sd289, 11'sd-963, 11'sd-595}},
{{12'sd1732, 13'sd-3178, 12'sd1510}, {12'sd1805, 6'sd-27, 10'sd-309}, {12'sd1531, 10'sd-473, 13'sd-3490}},
{{11'sd-911, 13'sd-2628, 13'sd-2838}, {13'sd4004, 13'sd-2660, 12'sd-1493}, {14'sd7875, 13'sd3453, 13'sd3284}},
{{9'sd245, 12'sd1499, 12'sd-1537}, {13'sd-2719, 10'sd-471, 10'sd-276}, {12'sd1370, 12'sd-1060, 8'sd-120}},
{{13'sd-2467, 12'sd1578, 12'sd-1352}, {10'sd-426, 9'sd-207, 11'sd-712}, {11'sd-771, 13'sd2870, 13'sd3146}},
{{12'sd-1176, 9'sd-134, 10'sd-351}, {12'sd-1850, 13'sd-2862, 13'sd-3093}, {12'sd-1603, 9'sd238, 10'sd464}},
{{10'sd468, 3'sd2, 13'sd-2185}, {12'sd1077, 13'sd2484, 12'sd1031}, {12'sd1541, 13'sd2156, 12'sd-1690}},
{{10'sd-504, 9'sd-207, 12'sd1505}, {13'sd3195, 12'sd1919, 13'sd-2823}, {13'sd2197, 12'sd1868, 13'sd-2660}},
{{12'sd-1085, 10'sd-429, 12'sd1099}, {12'sd-1971, 12'sd1382, 12'sd1101}, {10'sd-259, 13'sd-2295, 11'sd-673}},
{{12'sd1697, 13'sd3304, 12'sd-1115}, {12'sd-1082, 13'sd2627, 12'sd1368}, {13'sd2179, 12'sd1219, 11'sd-626}},
{{12'sd1245, 13'sd-2373, 12'sd1928}, {12'sd1945, 11'sd-998, 13'sd-2095}, {11'sd-943, 12'sd-1576, 11'sd974}},
{{13'sd-2454, 11'sd-641, 12'sd-1097}, {9'sd193, 10'sd-476, 12'sd-1497}, {11'sd-689, 12'sd-1823, 11'sd-654}},
{{11'sd-634, 7'sd-57, 12'sd1258}, {8'sd-109, 9'sd-187, 13'sd2823}, {8'sd-121, 11'sd729, 9'sd-185}},
{{9'sd247, 12'sd-1643, 10'sd290}, {11'sd-923, 7'sd60, 12'sd-1513}, {11'sd-861, 12'sd1549, 12'sd-1930}},
{{13'sd-2703, 12'sd-1550, 13'sd2154}, {11'sd851, 13'sd2075, 13'sd2500}, {10'sd-300, 9'sd225, 11'sd585}},
{{9'sd187, 13'sd2415, 13'sd2165}, {13'sd3025, 13'sd2996, 14'sd4517}, {10'sd317, 12'sd1481, 12'sd1735}},
{{13'sd2789, 13'sd-2673, 12'sd-1203}, {12'sd-1073, 12'sd-1191, 11'sd855}, {10'sd289, 12'sd-1589, 13'sd-2181}},
{{13'sd-3195, 12'sd-1539, 13'sd-3807}, {11'sd-611, 13'sd-3895, 8'sd93}, {11'sd-590, 10'sd281, 12'sd-1250}},
{{12'sd-1124, 12'sd-1657, 13'sd-2596}, {10'sd298, 9'sd200, 13'sd-3079}, {13'sd2226, 12'sd-1766, 12'sd1895}},
{{8'sd110, 12'sd1858, 13'sd2966}, {13'sd-2301, 12'sd-1140, 10'sd-392}, {12'sd1903, 9'sd-253, 11'sd-1001}},
{{13'sd3466, 10'sd-500, 13'sd-2309}, {13'sd2993, 13'sd-2098, 10'sd-390}, {13'sd3171, 9'sd-237, 12'sd-1122}},
{{11'sd929, 12'sd1292, 13'sd3077}, {13'sd-2419, 13'sd-2507, 9'sd159}, {12'sd-1201, 12'sd1134, 10'sd318}},
{{11'sd-597, 11'sd904, 12'sd-1030}, {13'sd2686, 12'sd-1892, 13'sd-3421}, {11'sd-733, 12'sd-1406, 9'sd139}}},
{
{{11'sd-577, 12'sd-1764, 12'sd-1375}, {11'sd-1008, 11'sd-590, 12'sd1281}, {13'sd2486, 11'sd-853, 13'sd2933}},
{{12'sd-1626, 12'sd1696, 12'sd-1263}, {13'sd2077, 13'sd2874, 11'sd650}, {12'sd1214, 11'sd874, 13'sd2228}},
{{13'sd3884, 12'sd1386, 12'sd-1437}, {12'sd1283, 11'sd-560, 12'sd1247}, {11'sd-945, 13'sd-3487, 13'sd-3126}},
{{9'sd-243, 10'sd317, 10'sd349}, {12'sd-1918, 8'sd-107, 11'sd-558}, {13'sd2749, 9'sd241, 12'sd1404}},
{{13'sd-2305, 11'sd810, 10'sd354}, {13'sd2372, 12'sd1068, 13'sd2745}, {11'sd923, 11'sd771, 11'sd1003}},
{{12'sd-1880, 12'sd1617, 13'sd-2119}, {12'sd1937, 12'sd1038, 13'sd2600}, {11'sd683, 12'sd1942, 11'sd-743}},
{{12'sd1532, 12'sd1070, 11'sd661}, {12'sd-1763, 11'sd-522, 12'sd1601}, {10'sd-476, 13'sd2191, 13'sd-2147}},
{{13'sd-2287, 12'sd-1996, 13'sd-2869}, {11'sd654, 12'sd1611, 9'sd-196}, {12'sd-1948, 13'sd2791, 12'sd1398}},
{{5'sd10, 12'sd1613, 12'sd1452}, {12'sd1333, 12'sd-1477, 8'sd78}, {10'sd489, 12'sd1899, 6'sd22}},
{{12'sd-1468, 11'sd-713, 12'sd-1136}, {11'sd-802, 11'sd715, 12'sd-1325}, {13'sd2087, 13'sd2313, 10'sd307}},
{{11'sd-918, 13'sd2154, 13'sd2363}, {13'sd2496, 13'sd3602, 10'sd428}, {11'sd-884, 12'sd-1895, 14'sd-4170}},
{{10'sd336, 12'sd-1643, 10'sd-486}, {12'sd1898, 13'sd-2067, 8'sd-70}, {9'sd135, 13'sd3573, 12'sd1819}},
{{12'sd1165, 9'sd242, 13'sd-2712}, {9'sd232, 14'sd-4200, 13'sd-3989}, {12'sd-1233, 13'sd-3460, 12'sd-1200}},
{{12'sd-1933, 11'sd621, 12'sd1347}, {11'sd724, 13'sd2379, 11'sd913}, {12'sd-1307, 13'sd-2108, 12'sd-1613}},
{{12'sd1698, 8'sd98, 11'sd-654}, {12'sd1889, 10'sd-312, 13'sd-2403}, {10'sd481, 12'sd-1492, 8'sd125}},
{{12'sd1465, 13'sd-3250, 12'sd-1891}, {9'sd226, 13'sd-2457, 10'sd-415}, {12'sd1047, 12'sd-1814, 13'sd2716}},
{{13'sd-2729, 12'sd-1321, 11'sd573}, {13'sd-2894, 13'sd-3817, 12'sd1895}, {13'sd-2347, 13'sd-2927, 12'sd-1900}},
{{13'sd-3027, 12'sd-1305, 14'sd-4529}, {12'sd1341, 13'sd3209, 14'sd-4311}, {12'sd-1244, 13'sd2070, 14'sd-4422}},
{{11'sd-868, 13'sd-3034, 13'sd-3067}, {11'sd764, 13'sd-2167, 13'sd-2424}, {8'sd-110, 11'sd-577, 12'sd-1781}},
{{12'sd1127, 13'sd-2454, 12'sd1042}, {10'sd-351, 12'sd-1187, 11'sd-553}, {9'sd209, 12'sd1604, 12'sd1074}},
{{12'sd1960, 12'sd1756, 10'sd506}, {12'sd-1896, 13'sd3081, 12'sd-1401}, {12'sd-1898, 10'sd259, 11'sd732}},
{{12'sd1500, 12'sd-1864, 13'sd3060}, {12'sd1416, 11'sd-968, 13'sd-2079}, {13'sd-2121, 10'sd477, 10'sd-419}},
{{13'sd3392, 13'sd2157, 13'sd2556}, {12'sd-1592, 12'sd-1667, 12'sd-1962}, {10'sd438, 9'sd173, 12'sd1840}},
{{10'sd474, 12'sd1315, 13'sd2766}, {12'sd1862, 12'sd1190, 8'sd101}, {12'sd1067, 12'sd1690, 13'sd2390}},
{{13'sd-2184, 11'sd554, 13'sd2700}, {13'sd2852, 12'sd1789, 14'sd4860}, {13'sd3220, 13'sd3077, 13'sd2198}},
{{10'sd342, 10'sd475, 12'sd1580}, {12'sd-1345, 12'sd1728, 10'sd-488}, {13'sd2484, 10'sd-307, 11'sd518}},
{{11'sd993, 13'sd-2441, 11'sd685}, {12'sd-1389, 12'sd-1939, 13'sd2238}, {12'sd-2040, 13'sd3129, 11'sd-941}},
{{12'sd-1057, 11'sd573, 9'sd236}, {12'sd-1342, 11'sd947, 12'sd-1831}, {11'sd676, 12'sd1417, 13'sd2135}},
{{12'sd1210, 13'sd2237, 12'sd1914}, {13'sd-3435, 12'sd1853, 13'sd-2896}, {10'sd-359, 13'sd-2704, 12'sd-1055}},
{{12'sd-1303, 12'sd1025, 12'sd-1124}, {13'sd-2145, 13'sd-3690, 9'sd239}, {11'sd603, 11'sd-772, 10'sd371}},
{{12'sd1639, 11'sd913, 10'sd-481}, {10'sd491, 13'sd-2063, 11'sd755}, {12'sd-1520, 13'sd-3162, 12'sd-1375}},
{{13'sd3075, 12'sd1675, 13'sd-2217}, {12'sd-1701, 12'sd-1216, 13'sd2828}, {11'sd-659, 13'sd2080, 12'sd1329}},
{{10'sd-451, 12'sd1761, 8'sd-119}, {10'sd-483, 13'sd2913, 12'sd-1643}, {12'sd1851, 13'sd2431, 13'sd-2451}},
{{9'sd-184, 10'sd297, 13'sd2248}, {12'sd1169, 12'sd1575, 12'sd-1975}, {13'sd-2714, 11'sd549, 13'sd-3467}},
{{8'sd-114, 8'sd-66, 13'sd2752}, {12'sd-1821, 12'sd-1896, 13'sd2506}, {12'sd1438, 8'sd103, 12'sd-1670}},
{{13'sd-3163, 12'sd1315, 13'sd-2656}, {8'sd105, 10'sd331, 12'sd1858}, {13'sd3024, 12'sd1577, 12'sd1814}},
{{13'sd3830, 12'sd-1877, 11'sd661}, {10'sd-280, 11'sd-709, 12'sd-1178}, {12'sd1304, 12'sd1045, 13'sd-2237}},
{{8'sd107, 13'sd-2735, 13'sd-3656}, {12'sd-1160, 13'sd-2457, 12'sd1194}, {13'sd2306, 11'sd701, 14'sd4240}},
{{12'sd-1104, 12'sd1621, 13'sd-2944}, {13'sd-2829, 10'sd350, 12'sd-1956}, {13'sd2747, 12'sd2045, 13'sd2164}},
{{13'sd-2245, 10'sd-262, 10'sd258}, {12'sd1724, 13'sd2120, 9'sd-205}, {13'sd-2706, 8'sd-65, 11'sd-568}},
{{11'sd-981, 11'sd900, 12'sd1805}, {13'sd2858, 12'sd1796, 13'sd2427}, {11'sd653, 10'sd505, 12'sd-2005}},
{{11'sd-867, 13'sd-2846, 11'sd-542}, {13'sd-2163, 13'sd2304, 8'sd-94}, {13'sd2733, 13'sd2807, 13'sd3709}},
{{11'sd825, 13'sd2780, 11'sd981}, {12'sd-1805, 12'sd1300, 13'sd2920}, {12'sd1144, 11'sd-971, 11'sd900}},
{{12'sd1146, 10'sd-397, 11'sd699}, {7'sd36, 9'sd-246, 11'sd-832}, {12'sd1994, 13'sd2650, 12'sd-1151}},
{{10'sd-400, 10'sd-487, 11'sd680}, {12'sd1617, 12'sd1275, 10'sd364}, {11'sd-563, 13'sd2285, 12'sd-1079}},
{{11'sd-1007, 10'sd-499, 10'sd-373}, {12'sd1675, 5'sd9, 13'sd2312}, {12'sd-1737, 11'sd626, 12'sd1458}},
{{12'sd1438, 9'sd-131, 11'sd611}, {13'sd-3048, 13'sd-3039, 11'sd975}, {12'sd-1553, 13'sd-2920, 11'sd-547}},
{{10'sd355, 11'sd582, 11'sd870}, {12'sd-1709, 13'sd2603, 11'sd-809}, {13'sd2490, 12'sd-1869, 7'sd-39}},
{{12'sd1866, 11'sd901, 13'sd-2434}, {12'sd-1943, 13'sd-2220, 13'sd-2340}, {12'sd-1522, 1'sd0, 13'sd2259}},
{{7'sd46, 11'sd649, 13'sd-2457}, {12'sd1630, 12'sd-1502, 11'sd-906}, {12'sd-1282, 9'sd224, 11'sd778}},
{{13'sd2157, 13'sd-2231, 12'sd1627}, {7'sd62, 10'sd-264, 11'sd826}, {12'sd-1306, 13'sd2557, 9'sd-191}},
{{8'sd112, 11'sd787, 13'sd-2856}, {12'sd-1833, 11'sd591, 11'sd733}, {13'sd-2920, 11'sd-938, 13'sd-2337}},
{{12'sd1181, 11'sd744, 13'sd-2048}, {12'sd-1146, 13'sd-2942, 13'sd-2281}, {12'sd1595, 11'sd874, 14'sd-4681}},
{{13'sd2392, 10'sd422, 11'sd886}, {13'sd2734, 13'sd-2603, 12'sd1522}, {12'sd-1138, 10'sd-389, 12'sd2012}},
{{13'sd2059, 12'sd-1108, 12'sd-1030}, {13'sd-2206, 13'sd-2305, 12'sd-1724}, {13'sd-2620, 12'sd-1251, 13'sd-3260}},
{{7'sd52, 12'sd1856, 11'sd-854}, {13'sd-2363, 13'sd-2286, 9'sd241}, {13'sd-2100, 13'sd-3030, 13'sd-3179}},
{{11'sd-643, 8'sd98, 12'sd1910}, {12'sd1478, 12'sd-1936, 11'sd-1008}, {12'sd-1324, 12'sd1512, 13'sd-2803}},
{{12'sd1955, 12'sd-1622, 12'sd1350}, {13'sd-2789, 13'sd2445, 12'sd1852}, {12'sd-1760, 11'sd-531, 12'sd1614}},
{{13'sd3094, 13'sd3959, 13'sd3448}, {12'sd1700, 13'sd-2166, 12'sd1212}, {12'sd1256, 12'sd1075, 13'sd2581}},
{{12'sd-1606, 13'sd2081, 13'sd2196}, {12'sd-1183, 9'sd-238, 12'sd1331}, {9'sd-207, 12'sd-1834, 12'sd1992}},
{{13'sd-2986, 11'sd-582, 11'sd861}, {12'sd-1279, 13'sd2260, 12'sd1196}, {13'sd-2268, 12'sd1071, 9'sd218}},
{{13'sd-2429, 10'sd-369, 13'sd-2303}, {13'sd-2594, 11'sd-764, 12'sd-1788}, {12'sd1497, 12'sd-2028, 13'sd2619}},
{{10'sd294, 12'sd-1401, 11'sd-938}, {13'sd2189, 13'sd-2165, 13'sd2061}, {13'sd2893, 13'sd2728, 9'sd131}},
{{10'sd364, 12'sd1616, 12'sd1040}, {10'sd462, 12'sd-1197, 12'sd1793}, {12'sd-1624, 12'sd1944, 11'sd867}}},
{
{{11'sd-557, 12'sd1854, 13'sd2479}, {12'sd1916, 12'sd-1344, 11'sd816}, {13'sd2093, 12'sd1199, 12'sd1083}},
{{13'sd2216, 11'sd585, 12'sd1359}, {10'sd-324, 11'sd-737, 13'sd-2413}, {12'sd-1725, 8'sd-116, 13'sd-2153}},
{{11'sd-897, 13'sd-2528, 13'sd-2344}, {12'sd-1891, 12'sd1817, 13'sd2117}, {8'sd118, 13'sd-3246, 11'sd-662}},
{{13'sd-2818, 13'sd2097, 13'sd2609}, {9'sd238, 12'sd-1983, 13'sd-2399}, {12'sd-1997, 11'sd673, 12'sd-2042}},
{{12'sd-1763, 12'sd1924, 13'sd2630}, {12'sd1112, 11'sd991, 13'sd2699}, {11'sd-821, 12'sd1809, 13'sd2736}},
{{11'sd839, 10'sd426, 13'sd2458}, {10'sd459, 12'sd-1185, 12'sd-1808}, {10'sd-329, 11'sd-767, 12'sd-1670}},
{{10'sd-471, 12'sd1617, 11'sd515}, {12'sd1055, 11'sd959, 12'sd-1502}, {12'sd-1479, 13'sd-3154, 8'sd70}},
{{11'sd895, 13'sd-2063, 13'sd-2498}, {11'sd-834, 10'sd380, 13'sd-2084}, {8'sd101, 13'sd-2228, 12'sd1442}},
{{11'sd-741, 11'sd597, 11'sd-728}, {10'sd-268, 11'sd943, 11'sd-599}, {12'sd-1669, 12'sd1388, 5'sd-10}},
{{11'sd-677, 12'sd-2008, 13'sd3141}, {13'sd-2131, 11'sd-974, 10'sd-302}, {13'sd-2850, 13'sd-3273, 11'sd-750}},
{{13'sd-3552, 11'sd-862, 12'sd1549}, {10'sd382, 12'sd1975, 12'sd-1158}, {10'sd-375, 12'sd1048, 12'sd2026}},
{{5'sd-8, 12'sd-1024, 9'sd234}, {12'sd1661, 11'sd-572, 7'sd-54}, {10'sd298, 12'sd1887, 12'sd1056}},
{{13'sd2618, 13'sd2320, 10'sd468}, {10'sd392, 10'sd346, 12'sd-1520}, {13'sd-3049, 9'sd224, 12'sd-1456}},
{{10'sd-333, 12'sd1560, 12'sd-1504}, {12'sd-1564, 11'sd-754, 10'sd-410}, {13'sd2585, 11'sd536, 13'sd-2448}},
{{12'sd-1158, 12'sd1806, 10'sd270}, {13'sd2715, 10'sd350, 12'sd1087}, {13'sd-2588, 9'sd-130, 13'sd2564}},
{{12'sd1318, 12'sd-1505, 10'sd-367}, {1'sd0, 13'sd2475, 9'sd180}, {12'sd-1544, 11'sd516, 12'sd1936}},
{{10'sd419, 11'sd-536, 12'sd-1060}, {13'sd2365, 6'sd-23, 11'sd699}, {12'sd1162, 11'sd587, 11'sd-856}},
{{12'sd-1831, 13'sd-3219, 13'sd-3335}, {13'sd-3263, 12'sd-1973, 12'sd1538}, {13'sd-3135, 9'sd253, 11'sd698}},
{{13'sd2278, 11'sd890, 12'sd1704}, {10'sd438, 13'sd-2579, 12'sd-1877}, {12'sd-1447, 11'sd-703, 10'sd-321}},
{{12'sd1449, 11'sd674, 11'sd-611}, {12'sd1333, 13'sd-2278, 12'sd2005}, {12'sd-1058, 9'sd221, 12'sd1566}},
{{11'sd877, 13'sd-3011, 11'sd983}, {12'sd-1482, 10'sd348, 11'sd628}, {12'sd-1307, 12'sd-1308, 12'sd1562}},
{{13'sd2473, 12'sd-1571, 12'sd-1500}, {13'sd3187, 13'sd2797, 9'sd-153}, {10'sd-299, 12'sd-1191, 9'sd-161}},
{{12'sd1471, 13'sd-2110, 12'sd-1814}, {12'sd-1561, 12'sd2017, 11'sd-846}, {11'sd736, 13'sd2924, 13'sd-2586}},
{{12'sd-2043, 13'sd2298, 12'sd-1493}, {12'sd-1742, 12'sd-1736, 12'sd1750}, {13'sd-3056, 12'sd-1179, 13'sd-2493}},
{{11'sd-620, 13'sd-3271, 10'sd-442}, {13'sd2169, 11'sd670, 11'sd-534}, {12'sd-1043, 12'sd1359, 12'sd1855}},
{{10'sd281, 11'sd988, 11'sd-1023}, {12'sd-1929, 13'sd-2068, 8'sd-75}, {11'sd679, 12'sd1497, 12'sd-1676}},
{{13'sd-2741, 10'sd283, 12'sd1059}, {11'sd634, 11'sd865, 12'sd-1402}, {13'sd2257, 12'sd-1630, 13'sd2628}},
{{10'sd498, 11'sd911, 12'sd-1137}, {10'sd-481, 12'sd-1484, 10'sd-501}, {9'sd-149, 13'sd-2480, 8'sd-121}},
{{12'sd-1126, 13'sd2363, 10'sd429}, {8'sd74, 12'sd1344, 11'sd633}, {12'sd-1070, 12'sd1840, 11'sd-851}},
{{12'sd-1061, 14'sd4192, 13'sd2595}, {13'sd-3072, 13'sd2665, 12'sd1293}, {13'sd-3021, 13'sd2301, 13'sd-2574}},
{{10'sd398, 13'sd2936, 7'sd47}, {12'sd-1703, 11'sd836, 13'sd-2146}, {12'sd-1653, 13'sd-2098, 9'sd160}},
{{7'sd-38, 12'sd1385, 12'sd-1298}, {12'sd-1392, 12'sd-1987, 11'sd-794}, {8'sd-83, 13'sd-2877, 11'sd870}},
{{11'sd970, 12'sd1787, 10'sd-393}, {12'sd1950, 12'sd1961, 13'sd2854}, {12'sd1386, 12'sd-1954, 13'sd2394}},
{{13'sd2553, 13'sd-2156, 7'sd-57}, {13'sd2535, 12'sd-1027, 11'sd-997}, {12'sd-1330, 9'sd163, 13'sd2054}},
{{13'sd-2245, 10'sd300, 13'sd2933}, {12'sd-1452, 12'sd1219, 12'sd1474}, {12'sd1764, 12'sd1613, 11'sd1009}},
{{12'sd-1343, 11'sd-630, 7'sd-55}, {12'sd-1433, 11'sd566, 13'sd-3062}, {13'sd2398, 8'sd-123, 13'sd2395}},
{{12'sd1797, 13'sd-3102, 12'sd-1238}, {11'sd598, 13'sd2625, 12'sd1220}, {12'sd-1841, 13'sd2668, 12'sd-1600}},
{{9'sd-225, 13'sd2636, 13'sd-2955}, {13'sd3805, 7'sd39, 13'sd-2414}, {12'sd1740, 13'sd3778, 13'sd-3175}},
{{12'sd-1129, 12'sd1165, 13'sd2345}, {12'sd-1862, 13'sd-2753, 12'sd2044}, {12'sd-1454, 11'sd791, 13'sd2552}},
{{12'sd-1408, 11'sd1012, 12'sd1908}, {11'sd-589, 11'sd-895, 11'sd578}, {12'sd-1127, 12'sd1117, 11'sd724}},
{{12'sd-1357, 10'sd-506, 13'sd2088}, {11'sd-731, 11'sd-926, 13'sd2554}, {13'sd2366, 12'sd-1296, 13'sd-2529}},
{{12'sd-1323, 11'sd-639, 12'sd1494}, {13'sd-2144, 12'sd2034, 13'sd-2728}, {12'sd-1215, 10'sd-282, 6'sd-26}},
{{11'sd678, 11'sd-970, 11'sd-697}, {12'sd1194, 13'sd-3352, 12'sd1544}, {10'sd-290, 12'sd-1793, 13'sd-2712}},
{{12'sd-1298, 13'sd-2909, 11'sd-835}, {13'sd2896, 12'sd1825, 12'sd-1517}, {13'sd2555, 12'sd1138, 12'sd-1954}},
{{12'sd-1725, 8'sd-86, 12'sd-1746}, {13'sd2746, 11'sd678, 12'sd1439}, {12'sd1160, 10'sd415, 12'sd-1255}},
{{11'sd981, 12'sd-1790, 11'sd-654}, {12'sd-1856, 12'sd-1269, 13'sd2723}, {13'sd3027, 13'sd2602, 6'sd-23}},
{{10'sd492, 11'sd645, 10'sd-276}, {10'sd-413, 12'sd-1511, 10'sd-462}, {13'sd-2571, 12'sd-1877, 13'sd-2299}},
{{11'sd-903, 9'sd-221, 12'sd2017}, {10'sd256, 13'sd2467, 13'sd2137}, {12'sd-1155, 11'sd-566, 13'sd2572}},
{{12'sd-1868, 10'sd-451, 9'sd-189}, {13'sd-2458, 12'sd-1881, 12'sd1185}, {12'sd1269, 10'sd-284, 8'sd-96}},
{{8'sd-117, 11'sd768, 12'sd1660}, {12'sd-1764, 11'sd-572, 13'sd2066}, {12'sd-1351, 11'sd-857, 13'sd2690}},
{{10'sd336, 13'sd-2292, 12'sd-1894}, {13'sd2858, 12'sd-1329, 12'sd1443}, {11'sd-873, 13'sd-2709, 13'sd-2086}},
{{12'sd-1236, 12'sd1340, 13'sd-2439}, {10'sd260, 12'sd1253, 11'sd720}, {12'sd1036, 13'sd-2365, 12'sd-1897}},
{{13'sd2111, 11'sd-804, 14'sd-4265}, {13'sd-2229, 13'sd2231, 13'sd-3717}, {13'sd-2206, 9'sd-218, 11'sd843}},
{{11'sd884, 13'sd2233, 12'sd-1992}, {10'sd466, 11'sd908, 9'sd-174}, {12'sd-1343, 13'sd-2640, 13'sd-2881}},
{{13'sd2769, 12'sd1306, 9'sd-158}, {13'sd3076, 11'sd-899, 8'sd105}, {10'sd432, 12'sd-1590, 12'sd-1226}},
{{13'sd2292, 11'sd-674, 11'sd842}, {13'sd2572, 5'sd-13, 12'sd1346}, {13'sd-2209, 12'sd1763, 12'sd-1204}},
{{11'sd-757, 11'sd-852, 13'sd-2911}, {13'sd3364, 13'sd3148, 13'sd-2075}, {13'sd2195, 12'sd1816, 12'sd1776}},
{{11'sd534, 9'sd175, 11'sd-845}, {12'sd-1917, 9'sd166, 7'sd41}, {13'sd2166, 13'sd-2064, 12'sd1972}},
{{13'sd-2133, 8'sd-106, 11'sd-562}, {13'sd-2182, 12'sd-1747, 13'sd2625}, {13'sd-3450, 10'sd-449, 13'sd-3163}},
{{13'sd-2119, 12'sd1923, 11'sd-542}, {12'sd-2042, 11'sd849, 12'sd1632}, {12'sd1057, 13'sd-2431, 13'sd2239}},
{{11'sd-842, 11'sd-708, 12'sd-1711}, {13'sd-2633, 13'sd-2501, 11'sd-972}, {12'sd1992, 11'sd792, 10'sd470}},
{{12'sd-1708, 12'sd1080, 13'sd2237}, {12'sd-1584, 11'sd823, 13'sd-2065}, {12'sd1400, 12'sd-1396, 12'sd-1063}},
{{12'sd1444, 10'sd274, 13'sd2758}, {12'sd1109, 13'sd-2590, 9'sd166}, {13'sd-2117, 11'sd-537, 13'sd2843}},
{{12'sd1272, 13'sd-2055, 9'sd-138}, {13'sd2363, 11'sd759, 12'sd1177}, {10'sd-437, 13'sd3580, 12'sd1384}}},
{
{{13'sd2337, 13'sd2445, 13'sd-2082}, {12'sd1151, 7'sd-44, 12'sd-1074}, {11'sd792, 5'sd10, 11'sd-1006}},
{{10'sd438, 12'sd1909, 9'sd176}, {11'sd951, 9'sd140, 13'sd2563}, {11'sd-581, 12'sd1231, 11'sd-875}},
{{12'sd-1522, 12'sd-1613, 11'sd818}, {12'sd1964, 11'sd-576, 12'sd-1312}, {13'sd2306, 11'sd-627, 13'sd3390}},
{{13'sd2314, 12'sd-1123, 12'sd1671}, {13'sd2938, 13'sd2323, 11'sd-675}, {11'sd873, 10'sd494, 12'sd-1175}},
{{13'sd2562, 10'sd-422, 10'sd-344}, {12'sd-1651, 13'sd3137, 13'sd-2175}, {13'sd2646, 11'sd-537, 13'sd3034}},
{{10'sd286, 12'sd-1155, 10'sd-265}, {12'sd-1088, 11'sd-630, 13'sd-2407}, {13'sd-2466, 12'sd1265, 12'sd1730}},
{{10'sd-388, 11'sd-564, 11'sd-515}, {10'sd421, 13'sd2120, 10'sd-372}, {11'sd955, 13'sd-2117, 10'sd-379}},
{{13'sd-3536, 9'sd-226, 13'sd-2285}, {12'sd-2035, 12'sd1397, 13'sd-2184}, {13'sd-2607, 12'sd-1703, 13'sd2224}},
{{12'sd-1911, 13'sd2750, 12'sd-1223}, {12'sd-1480, 9'sd229, 6'sd30}, {13'sd-2306, 11'sd-855, 8'sd91}},
{{6'sd-31, 12'sd2012, 11'sd873}, {12'sd1092, 12'sd1119, 13'sd2048}, {12'sd1629, 11'sd-1011, 11'sd1002}},
{{13'sd2665, 12'sd1730, 12'sd-1123}, {12'sd1881, 10'sd-508, 11'sd-681}, {13'sd-3382, 10'sd369, 13'sd-2474}},
{{11'sd875, 13'sd2580, 12'sd-1291}, {12'sd1591, 12'sd-1495, 13'sd2773}, {12'sd-1298, 12'sd1756, 11'sd814}},
{{13'sd-2954, 12'sd1657, 13'sd3279}, {11'sd979, 13'sd-2124, 10'sd509}, {13'sd-2583, 13'sd-2272, 13'sd-2289}},
{{13'sd-2217, 12'sd-1574, 11'sd-998}, {12'sd1601, 12'sd1611, 13'sd2285}, {9'sd-175, 10'sd429, 9'sd224}},
{{12'sd-1391, 9'sd143, 13'sd-2680}, {12'sd1560, 12'sd1300, 9'sd243}, {12'sd-1817, 11'sd669, 13'sd-2484}},
{{11'sd1017, 10'sd509, 13'sd2071}, {11'sd995, 12'sd1393, 13'sd2524}, {12'sd-1564, 12'sd1639, 11'sd-779}},
{{9'sd215, 8'sd96, 13'sd2783}, {12'sd-1133, 12'sd-1623, 13'sd2337}, {13'sd-2548, 12'sd1335, 11'sd993}},
{{14'sd-5406, 12'sd1047, 12'sd-2031}, {13'sd-3046, 12'sd-1948, 9'sd-172}, {13'sd3774, 13'sd2984, 13'sd2139}},
{{11'sd844, 12'sd1933, 13'sd2434}, {12'sd1314, 8'sd-117, 13'sd2259}, {11'sd-948, 11'sd623, 9'sd-167}},
{{11'sd-651, 13'sd-2810, 12'sd-1600}, {11'sd529, 12'sd1322, 12'sd1756}, {9'sd-253, 12'sd-1427, 12'sd-1863}},
{{12'sd1122, 12'sd-1265, 11'sd-595}, {13'sd2590, 11'sd-751, 13'sd-2187}, {11'sd-566, 11'sd939, 12'sd1169}},
{{12'sd-1624, 9'sd246, 12'sd1811}, {9'sd-213, 12'sd1470, 13'sd-2490}, {13'sd-2759, 8'sd107, 12'sd-1802}},
{{11'sd867, 8'sd-68, 12'sd-1824}, {12'sd-1109, 13'sd-2855, 11'sd-794}, {12'sd1133, 13'sd-2235, 10'sd-506}},
{{13'sd2789, 11'sd-1022, 13'sd2101}, {13'sd2072, 9'sd-199, 12'sd-1916}, {13'sd-2271, 12'sd-1691, 12'sd-1605}},
{{13'sd-2390, 11'sd995, 2'sd-1}, {11'sd985, 11'sd-811, 13'sd3895}, {6'sd27, 13'sd3277, 14'sd4339}},
{{9'sd-153, 13'sd-2387, 6'sd-18}, {12'sd-1024, 10'sd510, 11'sd792}, {13'sd-2206, 12'sd-1249, 7'sd-36}},
{{12'sd-1232, 12'sd1838, 12'sd-1177}, {12'sd-1598, 13'sd2197, 13'sd2207}, {11'sd-868, 12'sd2011, 13'sd2934}},
{{13'sd-2890, 11'sd-796, 12'sd-1936}, {11'sd-998, 12'sd1230, 10'sd-486}, {12'sd-1075, 12'sd1830, 9'sd128}},
{{9'sd-230, 9'sd187, 10'sd-506}, {9'sd130, 12'sd1281, 13'sd2192}, {10'sd-307, 12'sd1126, 9'sd-207}},
{{6'sd17, 11'sd-660, 8'sd-86}, {12'sd-1489, 7'sd53, 12'sd-1403}, {13'sd-2230, 10'sd330, 11'sd998}},
{{11'sd-838, 13'sd2342, 12'sd-1096}, {11'sd-749, 11'sd599, 12'sd-2035}, {12'sd1885, 9'sd-163, 10'sd-489}},
{{12'sd1551, 12'sd-1082, 11'sd-637}, {12'sd1478, 12'sd-1731, 12'sd-1678}, {12'sd-1158, 12'sd1928, 12'sd-1888}},
{{13'sd2275, 12'sd1416, 13'sd2742}, {7'sd-48, 12'sd1408, 11'sd864}, {10'sd-348, 12'sd-1410, 12'sd-1925}},
{{12'sd1959, 11'sd-614, 12'sd-1643}, {13'sd-2558, 12'sd1549, 13'sd-2224}, {13'sd2308, 12'sd-1125, 11'sd-709}},
{{11'sd-1006, 13'sd2556, 13'sd2133}, {12'sd1921, 11'sd673, 12'sd-1383}, {9'sd-203, 9'sd-161, 12'sd-1782}},
{{11'sd-923, 13'sd2459, 7'sd-37}, {13'sd2507, 12'sd-1370, 12'sd-1128}, {12'sd-1120, 12'sd-1528, 13'sd2159}},
{{11'sd-584, 12'sd-1856, 13'sd-2339}, {11'sd756, 12'sd1798, 9'sd-239}, {12'sd1234, 9'sd136, 13'sd2748}},
{{13'sd2509, 12'sd-1131, 12'sd1428}, {12'sd1037, 12'sd1136, 9'sd-177}, {11'sd850, 10'sd-258, 12'sd1453}},
{{13'sd-2183, 11'sd813, 12'sd1698}, {10'sd475, 12'sd-1681, 12'sd1569}, {11'sd-798, 12'sd-1319, 8'sd-98}},
{{9'sd-129, 10'sd-348, 13'sd-3251}, {13'sd2133, 11'sd-809, 12'sd1032}, {13'sd2793, 12'sd-1420, 12'sd1966}},
{{11'sd-857, 11'sd900, 8'sd96}, {12'sd-1166, 13'sd-2193, 13'sd-2252}, {11'sd580, 12'sd1255, 12'sd1368}},
{{12'sd1421, 13'sd2317, 10'sd-301}, {12'sd2037, 12'sd-1681, 9'sd205}, {13'sd-2352, 12'sd-1607, 13'sd2916}},
{{11'sd-719, 7'sd59, 12'sd-2030}, {12'sd1328, 12'sd-1133, 13'sd2546}, {12'sd2001, 13'sd-2242, 12'sd1207}},
{{12'sd1719, 9'sd-214, 12'sd-2047}, {12'sd-1457, 13'sd-2746, 11'sd549}, {13'sd-2997, 11'sd535, 13'sd-2251}},
{{11'sd-654, 12'sd1081, 11'sd704}, {11'sd-893, 10'sd463, 13'sd-2265}, {13'sd-2094, 8'sd-119, 9'sd-237}},
{{8'sd68, 13'sd-2145, 7'sd40}, {12'sd-1342, 11'sd820, 13'sd2212}, {12'sd1081, 10'sd342, 13'sd2844}},
{{11'sd-550, 11'sd578, 12'sd1512}, {13'sd-2486, 12'sd1939, 11'sd-625}, {12'sd-1681, 13'sd2552, 11'sd-665}},
{{12'sd2039, 12'sd1768, 10'sd424}, {11'sd-915, 12'sd1883, 11'sd718}, {12'sd1125, 10'sd-274, 12'sd-1484}},
{{12'sd1280, 13'sd2481, 12'sd1823}, {12'sd-1075, 13'sd2473, 13'sd-2549}, {12'sd1302, 11'sd-761, 13'sd-2856}},
{{9'sd-226, 12'sd1084, 13'sd2155}, {9'sd128, 13'sd-2202, 10'sd-453}, {12'sd1150, 13'sd2425, 11'sd670}},
{{12'sd-1434, 11'sd788, 11'sd805}, {11'sd1021, 10'sd397, 10'sd-261}, {12'sd1876, 7'sd36, 13'sd-2547}},
{{11'sd-716, 13'sd-2536, 13'sd-2219}, {12'sd-1633, 13'sd-2512, 10'sd-334}, {10'sd427, 9'sd235, 12'sd-1668}},
{{12'sd-1589, 12'sd-1896, 12'sd1213}, {10'sd-502, 12'sd-2045, 13'sd-2570}, {14'sd4288, 12'sd-1216, 13'sd3276}},
{{12'sd-1138, 11'sd-974, 13'sd-2309}, {12'sd-1963, 11'sd925, 9'sd-215}, {11'sd-980, 12'sd1785, 13'sd2630}},
{{11'sd-1000, 11'sd-568, 13'sd-2676}, {13'sd-2281, 12'sd-1297, 13'sd-2180}, {9'sd-235, 12'sd-1755, 13'sd-2517}},
{{13'sd-2179, 13'sd2144, 12'sd1548}, {13'sd-2272, 13'sd-2658, 10'sd-399}, {11'sd889, 10'sd-390, 13'sd-2478}},
{{11'sd862, 9'sd-162, 12'sd-1566}, {11'sd-961, 13'sd-2083, 12'sd-1250}, {12'sd1371, 10'sd-455, 12'sd1045}},
{{13'sd-2785, 13'sd-3474, 8'sd-86}, {12'sd-1371, 10'sd305, 11'sd923}, {12'sd1967, 10'sd-360, 10'sd-481}},
{{12'sd-1950, 10'sd-411, 12'sd1133}, {11'sd942, 12'sd-1250, 13'sd-2208}, {10'sd414, 12'sd-1175, 13'sd2478}},
{{13'sd-2355, 12'sd-1451, 12'sd2020}, {11'sd701, 12'sd-2030, 12'sd-1261}, {12'sd2002, 13'sd2492, 11'sd-603}},
{{12'sd-1032, 9'sd221, 12'sd-1265}, {12'sd-1982, 13'sd2253, 13'sd2104}, {13'sd-2294, 13'sd2578, 13'sd2718}},
{{11'sd-606, 13'sd-2558, 13'sd-2569}, {10'sd-377, 13'sd2213, 11'sd938}, {10'sd483, 11'sd-875, 11'sd-793}},
{{10'sd-487, 12'sd-1164, 11'sd-768}, {13'sd2345, 12'sd1135, 11'sd-858}, {12'sd-1170, 9'sd-190, 13'sd2860}},
{{9'sd-229, 10'sd428, 10'sd-468}, {11'sd-551, 12'sd1751, 13'sd-2953}, {10'sd489, 12'sd-1663, 13'sd-2738}}},
{
{{13'sd-2961, 13'sd-3627, 13'sd-2775}, {12'sd-1218, 12'sd-1598, 10'sd-299}, {13'sd2326, 10'sd507, 13'sd3244}},
{{12'sd1290, 12'sd-1472, 13'sd2113}, {9'sd-193, 13'sd2266, 13'sd3877}, {12'sd-1249, 12'sd1599, 13'sd-2323}},
{{12'sd1416, 13'sd-2408, 10'sd368}, {12'sd1709, 12'sd-1211, 13'sd2253}, {12'sd1225, 11'sd-601, 11'sd-977}},
{{12'sd1532, 13'sd-2309, 10'sd-414}, {12'sd-1504, 12'sd1460, 12'sd1412}, {12'sd1360, 12'sd1781, 13'sd3148}},
{{12'sd-1670, 12'sd1585, 9'sd223}, {11'sd839, 12'sd1092, 11'sd784}, {12'sd-1821, 12'sd-1322, 10'sd-265}},
{{12'sd1378, 10'sd480, 11'sd-657}, {11'sd-928, 9'sd-218, 11'sd657}, {11'sd-866, 11'sd826, 10'sd490}},
{{8'sd-74, 12'sd1174, 13'sd2389}, {9'sd-173, 13'sd-2567, 12'sd-2020}, {11'sd-667, 13'sd-3230, 12'sd-1292}},
{{14'sd-4282, 12'sd-1753, 10'sd-261}, {11'sd827, 7'sd-38, 13'sd-2560}, {13'sd2916, 13'sd2683, 12'sd-1427}},
{{13'sd3166, 13'sd2899, 11'sd-738}, {12'sd1418, 12'sd-1419, 13'sd2093}, {13'sd2773, 10'sd-376, 13'sd-2061}},
{{11'sd-727, 9'sd170, 13'sd2251}, {13'sd-3844, 12'sd-1881, 11'sd-614}, {13'sd-3035, 10'sd-395, 11'sd-702}},
{{10'sd-492, 13'sd3351, 8'sd-94}, {14'sd-4232, 12'sd-1737, 12'sd-1880}, {12'sd1628, 12'sd1171, 13'sd2277}},
{{12'sd1245, 12'sd1965, 13'sd2656}, {12'sd1199, 12'sd2031, 12'sd1388}, {12'sd1949, 10'sd-338, 11'sd-517}},
{{13'sd-3177, 11'sd-642, 13'sd-2082}, {11'sd-974, 12'sd-1815, 10'sd-427}, {10'sd464, 13'sd-2289, 12'sd1027}},
{{11'sd-753, 13'sd2417, 11'sd807}, {12'sd-1646, 13'sd-2578, 11'sd-650}, {13'sd2811, 13'sd-2337, 11'sd854}},
{{12'sd-1283, 12'sd-1311, 12'sd-1571}, {12'sd-1083, 11'sd-1012, 12'sd1091}, {13'sd-2424, 12'sd1210, 13'sd-2341}},
{{10'sd294, 12'sd-1232, 11'sd-948}, {12'sd-1971, 7'sd34, 11'sd813}, {11'sd-551, 13'sd2824, 10'sd400}},
{{11'sd883, 12'sd1433, 12'sd-1053}, {12'sd-1322, 12'sd-1277, 13'sd2928}, {13'sd-2298, 13'sd-2601, 10'sd439}},
{{13'sd-2830, 11'sd981, 12'sd-1258}, {13'sd-2220, 13'sd2944, 13'sd2119}, {13'sd-3426, 13'sd-2938, 14'sd-4883}},
{{9'sd-171, 12'sd1994, 12'sd1429}, {9'sd-213, 11'sd594, 4'sd5}, {13'sd2223, 9'sd176, 12'sd1497}},
{{12'sd-1092, 12'sd1618, 12'sd1564}, {10'sd492, 12'sd1148, 12'sd-1754}, {12'sd-1870, 13'sd-2108, 13'sd3079}},
{{12'sd1354, 13'sd2638, 13'sd2608}, {11'sd715, 13'sd2157, 9'sd-239}, {13'sd2677, 13'sd-2514, 9'sd-147}},
{{9'sd226, 12'sd-1555, 13'sd2208}, {12'sd1688, 12'sd-1765, 9'sd159}, {13'sd-2537, 12'sd-1181, 11'sd-769}},
{{10'sd-263, 13'sd2256, 12'sd-1241}, {13'sd2530, 10'sd-321, 13'sd2274}, {12'sd-1840, 12'sd-1236, 12'sd1459}},
{{12'sd1078, 10'sd-357, 11'sd685}, {13'sd-3040, 13'sd2415, 10'sd353}, {12'sd-1751, 12'sd1530, 13'sd-2193}},
{{13'sd2975, 13'sd-2740, 12'sd1364}, {13'sd3779, 12'sd1397, 12'sd-1277}, {11'sd-961, 13'sd-2210, 11'sd-548}},
{{12'sd1684, 7'sd44, 12'sd1413}, {7'sd56, 12'sd-1095, 13'sd2522}, {8'sd69, 11'sd-697, 13'sd-2331}},
{{12'sd-1077, 13'sd-2158, 12'sd1185}, {11'sd814, 13'sd-2276, 10'sd-412}, {13'sd2100, 13'sd2361, 13'sd-2059}},
{{12'sd1352, 12'sd-1952, 8'sd73}, {12'sd1799, 12'sd1297, 11'sd-593}, {9'sd-253, 12'sd1147, 13'sd2287}},
{{12'sd1605, 13'sd2427, 12'sd1956}, {13'sd-2236, 12'sd-1146, 12'sd-1322}, {12'sd-1899, 12'sd-1905, 9'sd-222}},
{{12'sd-1860, 11'sd-1019, 12'sd1381}, {12'sd1453, 12'sd-1031, 11'sd-598}, {11'sd816, 11'sd-565, 13'sd-2495}},
{{13'sd2706, 13'sd2224, 10'sd505}, {13'sd3090, 11'sd965, 10'sd-347}, {11'sd-518, 13'sd2691, 12'sd-1111}},
{{13'sd-2105, 12'sd1959, 13'sd-3256}, {12'sd1510, 10'sd-288, 10'sd-316}, {12'sd1458, 13'sd-2633, 11'sd-763}},
{{12'sd-1924, 12'sd1591, 13'sd2541}, {13'sd2229, 12'sd-1613, 11'sd-554}, {10'sd433, 12'sd1070, 12'sd1764}},
{{11'sd892, 8'sd-95, 12'sd-1194}, {11'sd694, 10'sd406, 9'sd133}, {11'sd-971, 12'sd1355, 13'sd-2900}},
{{12'sd1132, 10'sd-367, 12'sd-1949}, {10'sd300, 13'sd-2729, 11'sd-982}, {12'sd-1557, 12'sd-1307, 13'sd2378}},
{{13'sd2642, 13'sd-2645, 12'sd1970}, {8'sd-117, 13'sd-2108, 12'sd-1076}, {12'sd1524, 7'sd-36, 11'sd-726}},
{{11'sd549, 12'sd1456, 10'sd433}, {13'sd-2269, 12'sd1681, 13'sd2088}, {10'sd-317, 13'sd2208, 12'sd1821}},
{{11'sd569, 13'sd2331, 9'sd-180}, {12'sd1777, 13'sd-2677, 12'sd-1303}, {13'sd-3374, 12'sd1776, 12'sd1584}},
{{13'sd-3490, 8'sd-92, 13'sd-2700}, {11'sd-956, 12'sd1315, 13'sd3467}, {12'sd-1909, 13'sd2232, 12'sd2032}},
{{8'sd70, 12'sd-1995, 12'sd1809}, {12'sd1185, 12'sd1724, 12'sd-1300}, {7'sd50, 11'sd691, 13'sd-2112}},
{{9'sd168, 10'sd401, 12'sd1852}, {12'sd1478, 12'sd1704, 12'sd-1498}, {13'sd3191, 12'sd1363, 12'sd2022}},
{{11'sd-794, 11'sd-866, 8'sd-91}, {12'sd-1704, 9'sd-135, 11'sd945}, {13'sd2500, 13'sd2068, 12'sd1713}},
{{13'sd-2475, 12'sd1959, 8'sd127}, {12'sd-1516, 12'sd-1781, 13'sd2870}, {13'sd2115, 13'sd2772, 13'sd2048}},
{{11'sd-576, 13'sd2071, 12'sd1780}, {13'sd2572, 11'sd669, 10'sd-350}, {13'sd2230, 13'sd2104, 11'sd-647}},
{{11'sd-1011, 8'sd-100, 11'sd599}, {13'sd-2906, 12'sd-1913, 12'sd-1543}, {12'sd2019, 11'sd767, 12'sd-1350}},
{{8'sd-120, 12'sd1847, 11'sd-993}, {11'sd-853, 12'sd1074, 12'sd1162}, {13'sd-2587, 12'sd-1649, 12'sd1857}},
{{10'sd-483, 12'sd1647, 10'sd-406}, {13'sd2395, 13'sd-2540, 10'sd318}, {10'sd-368, 13'sd-2506, 13'sd3126}},
{{13'sd3213, 12'sd1980, 9'sd-167}, {12'sd1394, 9'sd-193, 10'sd276}, {11'sd643, 12'sd-1240, 12'sd-1841}},
{{12'sd1638, 11'sd738, 12'sd-1962}, {10'sd302, 12'sd-1486, 12'sd1151}, {12'sd-1558, 13'sd2460, 12'sd1177}},
{{13'sd2500, 7'sd-47, 9'sd-132}, {12'sd-1577, 10'sd-510, 13'sd-2129}, {12'sd1573, 13'sd-2065, 9'sd234}},
{{10'sd467, 9'sd196, 8'sd73}, {12'sd1672, 12'sd-1910, 11'sd793}, {13'sd2460, 11'sd-836, 13'sd2092}},
{{11'sd602, 12'sd-1160, 12'sd-1198}, {11'sd887, 13'sd-2147, 10'sd474}, {11'sd761, 12'sd-1076, 13'sd-2584}},
{{13'sd3965, 13'sd3514, 11'sd871}, {13'sd2148, 11'sd685, 12'sd-1879}, {14'sd-4997, 13'sd-3218, 10'sd287}},
{{11'sd-905, 12'sd-1658, 12'sd-1276}, {9'sd-186, 9'sd172, 10'sd-493}, {12'sd-1581, 12'sd1129, 9'sd-230}},
{{11'sd585, 12'sd-1298, 12'sd2004}, {9'sd-223, 13'sd2400, 12'sd1664}, {13'sd2052, 12'sd1509, 12'sd-1367}},
{{11'sd755, 12'sd1242, 13'sd-2146}, {9'sd191, 11'sd-879, 12'sd1804}, {11'sd-995, 9'sd-215, 12'sd-1775}},
{{11'sd623, 11'sd972, 13'sd-2144}, {13'sd3040, 13'sd2409, 12'sd-1828}, {12'sd1177, 12'sd1239, 11'sd879}},
{{9'sd-225, 12'sd1126, 13'sd-2232}, {12'sd-1503, 12'sd1412, 13'sd-2696}, {6'sd28, 13'sd-2882, 12'sd1452}},
{{14'sd-4116, 13'sd-2428, 12'sd1142}, {13'sd-3378, 12'sd1826, 11'sd-983}, {12'sd-1354, 12'sd1778, 11'sd-732}},
{{12'sd-1923, 13'sd-2701, 12'sd1154}, {13'sd2571, 13'sd2171, 10'sd367}, {11'sd731, 12'sd-2016, 13'sd2770}},
{{12'sd1106, 10'sd-308, 12'sd-1506}, {12'sd1388, 13'sd-2262, 12'sd1432}, {10'sd-409, 13'sd-2433, 10'sd-419}},
{{13'sd-2660, 13'sd-2462, 13'sd2122}, {12'sd1403, 12'sd1740, 13'sd2574}, {13'sd3230, 9'sd-224, 12'sd1783}},
{{13'sd2491, 12'sd-1555, 12'sd1856}, {11'sd550, 10'sd-266, 12'sd-1677}, {11'sd846, 11'sd-741, 12'sd1212}},
{{12'sd1831, 10'sd-267, 12'sd-1673}, {12'sd1058, 11'sd-550, 13'sd2968}, {9'sd135, 12'sd1469, 12'sd1176}}},
{
{{8'sd121, 13'sd-2730, 12'sd1685}, {12'sd1287, 10'sd-287, 11'sd-701}, {13'sd2062, 12'sd-1462, 10'sd497}},
{{12'sd-1920, 13'sd-2609, 13'sd-2162}, {12'sd-1887, 10'sd-440, 11'sd-753}, {13'sd-2068, 10'sd-499, 12'sd1756}},
{{13'sd-3408, 10'sd458, 12'sd1067}, {12'sd-1582, 13'sd2652, 11'sd-927}, {12'sd1317, 11'sd-660, 12'sd2047}},
{{11'sd569, 12'sd1463, 9'sd146}, {12'sd2022, 10'sd258, 12'sd1926}, {12'sd1034, 12'sd-1366, 12'sd1135}},
{{13'sd-2628, 12'sd-1236, 12'sd-1806}, {12'sd1321, 12'sd-1791, 10'sd-284}, {12'sd-1047, 9'sd-139, 13'sd2126}},
{{8'sd65, 13'sd-2094, 8'sd77}, {11'sd-1003, 13'sd2134, 8'sd-118}, {13'sd2186, 12'sd-1612, 11'sd567}},
{{12'sd-1481, 11'sd711, 12'sd-1412}, {12'sd1173, 10'sd395, 12'sd1362}, {11'sd-942, 10'sd-391, 13'sd2152}},
{{13'sd-2951, 12'sd-1820, 12'sd1804}, {7'sd46, 8'sd69, 12'sd1621}, {13'sd-3234, 13'sd-2117, 5'sd-13}},
{{12'sd-1385, 10'sd388, 12'sd-1975}, {12'sd1060, 12'sd-1660, 13'sd2455}, {11'sd795, 11'sd-584, 12'sd-1847}},
{{13'sd2076, 13'sd-2923, 13'sd2590}, {12'sd-1415, 12'sd1242, 11'sd676}, {12'sd1462, 13'sd2279, 13'sd-2869}},
{{13'sd2979, 13'sd-2348, 11'sd733}, {12'sd1907, 12'sd-1358, 10'sd299}, {10'sd-496, 13'sd2226, 12'sd-1134}},
{{10'sd-367, 11'sd-756, 12'sd-1228}, {13'sd2164, 12'sd1461, 12'sd-1075}, {12'sd1062, 11'sd785, 13'sd-2625}},
{{5'sd15, 10'sd490, 10'sd-448}, {9'sd176, 13'sd2271, 9'sd-134}, {12'sd1223, 5'sd-15, 12'sd1221}},
{{12'sd-1067, 11'sd514, 13'sd-2801}, {10'sd442, 13'sd-2552, 11'sd-714}, {13'sd2098, 13'sd2337, 12'sd1817}},
{{11'sd-792, 11'sd897, 11'sd625}, {11'sd-574, 11'sd-954, 13'sd-2115}, {12'sd-1580, 11'sd-703, 11'sd919}},
{{8'sd-100, 10'sd329, 12'sd1049}, {13'sd-2615, 12'sd-1911, 11'sd923}, {13'sd-3121, 13'sd-2704, 12'sd1106}},
{{12'sd1758, 10'sd-407, 13'sd-2123}, {13'sd2412, 13'sd2182, 12'sd-1727}, {12'sd-1882, 11'sd810, 12'sd1222}},
{{13'sd-2538, 11'sd703, 12'sd1203}, {8'sd85, 12'sd2039, 12'sd1464}, {12'sd-1646, 12'sd1090, 11'sd798}},
{{13'sd-2232, 13'sd-2082, 11'sd740}, {12'sd1322, 12'sd-1064, 11'sd841}, {11'sd-698, 13'sd-2055, 13'sd2554}},
{{12'sd-1032, 11'sd831, 11'sd685}, {12'sd-1770, 8'sd86, 12'sd1375}, {11'sd-838, 13'sd-3128, 9'sd181}},
{{13'sd2722, 13'sd2492, 11'sd-859}, {12'sd1107, 12'sd1226, 11'sd-705}, {11'sd744, 12'sd-1908, 9'sd-246}},
{{13'sd3005, 11'sd-759, 12'sd1878}, {11'sd-775, 13'sd2579, 12'sd1260}, {13'sd-2260, 13'sd3058, 11'sd-943}},
{{12'sd-1815, 13'sd-2531, 12'sd-1170}, {8'sd-71, 13'sd-2395, 12'sd-1874}, {13'sd-2551, 12'sd-1054, 10'sd310}},
{{12'sd-1228, 13'sd2344, 7'sd38}, {11'sd-546, 13'sd-2674, 12'sd-1688}, {11'sd-719, 11'sd-863, 12'sd-1268}},
{{12'sd1423, 9'sd-219, 10'sd-391}, {12'sd-1738, 12'sd1184, 13'sd2218}, {11'sd-961, 13'sd3672, 13'sd2595}},
{{11'sd768, 11'sd865, 10'sd358}, {12'sd1842, 11'sd795, 12'sd-1413}, {11'sd-867, 9'sd206, 11'sd-958}},
{{11'sd733, 8'sd-76, 9'sd-208}, {12'sd1967, 12'sd1452, 7'sd-62}, {13'sd2815, 10'sd391, 13'sd2621}},
{{12'sd1960, 9'sd174, 11'sd730}, {13'sd-2507, 11'sd673, 13'sd2275}, {13'sd-2245, 12'sd1617, 12'sd-1091}},
{{8'sd-109, 10'sd-309, 12'sd-1735}, {12'sd1091, 12'sd-1107, 12'sd1811}, {10'sd451, 13'sd2475, 12'sd-1819}},
{{12'sd1954, 12'sd1295, 13'sd-2764}, {12'sd1230, 13'sd2050, 10'sd402}, {12'sd1119, 13'sd2254, 12'sd-1579}},
{{10'sd262, 12'sd-1481, 11'sd-775}, {13'sd2443, 12'sd-1811, 12'sd1024}, {10'sd504, 12'sd-1932, 11'sd-1016}},
{{10'sd365, 11'sd993, 12'sd-1281}, {9'sd-177, 11'sd-681, 13'sd2242}, {12'sd-1296, 11'sd-664, 11'sd-790}},
{{12'sd-1366, 11'sd767, 12'sd1190}, {13'sd-2538, 11'sd-676, 13'sd-2728}, {11'sd623, 13'sd2491, 13'sd-2618}},
{{12'sd1978, 13'sd2385, 13'sd2417}, {11'sd867, 12'sd-1553, 12'sd-1805}, {12'sd-1526, 7'sd61, 11'sd949}},
{{13'sd2339, 12'sd1330, 12'sd-2044}, {12'sd1047, 10'sd-395, 12'sd-1354}, {13'sd-2511, 9'sd-169, 7'sd-40}},
{{9'sd-181, 12'sd-1625, 12'sd-1192}, {9'sd198, 12'sd-1229, 11'sd969}, {12'sd1398, 12'sd-1438, 13'sd2290}},
{{13'sd2470, 12'sd-1118, 7'sd-46}, {13'sd-2605, 11'sd-848, 12'sd-1853}, {13'sd-2523, 7'sd60, 12'sd-1236}},
{{10'sd-394, 11'sd782, 12'sd-1877}, {11'sd642, 12'sd1920, 12'sd1674}, {10'sd-409, 13'sd3019, 10'sd488}},
{{9'sd-250, 13'sd-2213, 13'sd-2073}, {11'sd-702, 12'sd1572, 11'sd948}, {12'sd-1429, 13'sd-2494, 11'sd-681}},
{{13'sd-2663, 12'sd-1195, 13'sd2364}, {11'sd782, 11'sd685, 12'sd1580}, {12'sd-2032, 10'sd-488, 12'sd-1124}},
{{13'sd2335, 13'sd2674, 12'sd1524}, {11'sd-1006, 10'sd-275, 12'sd1731}, {12'sd-1378, 11'sd-812, 13'sd-2074}},
{{10'sd-356, 12'sd1871, 12'sd-1828}, {11'sd-514, 12'sd-1927, 12'sd-1089}, {13'sd2506, 12'sd-1654, 13'sd2295}},
{{11'sd-552, 12'sd-1419, 10'sd-256}, {11'sd961, 11'sd606, 13'sd-2410}, {9'sd-194, 12'sd-1398, 12'sd1300}},
{{12'sd1823, 12'sd-1519, 9'sd-204}, {12'sd1823, 13'sd2162, 11'sd647}, {13'sd2803, 11'sd945, 11'sd1003}},
{{13'sd2150, 12'sd-1751, 13'sd2294}, {10'sd348, 11'sd-852, 10'sd-340}, {12'sd-1678, 12'sd1757, 10'sd-478}},
{{10'sd504, 12'sd-1777, 13'sd2178}, {13'sd-2337, 6'sd-20, 13'sd-2124}, {13'sd2096, 12'sd1189, 13'sd3343}},
{{8'sd109, 13'sd2162, 12'sd-1743}, {11'sd-1009, 12'sd1851, 11'sd795}, {10'sd271, 13'sd2434, 13'sd-2941}},
{{12'sd1084, 11'sd-814, 8'sd-67}, {13'sd-2460, 12'sd1401, 13'sd-2291}, {12'sd-1777, 11'sd-715, 13'sd-2150}},
{{12'sd-1323, 13'sd2228, 12'sd1936}, {11'sd775, 10'sd269, 12'sd-1642}, {11'sd-905, 12'sd1983, 12'sd1667}},
{{11'sd729, 13'sd-2273, 13'sd2373}, {12'sd-1985, 11'sd-612, 12'sd1449}, {12'sd-1314, 11'sd-582, 9'sd-135}},
{{12'sd1787, 12'sd-1088, 12'sd-1378}, {12'sd-1705, 11'sd-593, 11'sd1007}, {11'sd575, 11'sd-516, 12'sd1628}},
{{11'sd628, 13'sd-2729, 12'sd-1512}, {11'sd-765, 12'sd-1312, 11'sd672}, {10'sd-417, 12'sd1586, 12'sd-1512}},
{{12'sd-1196, 11'sd-853, 10'sd-459}, {13'sd2214, 12'sd-1935, 9'sd247}, {13'sd2667, 12'sd1150, 13'sd2355}},
{{11'sd874, 12'sd1735, 12'sd1933}, {12'sd-1941, 12'sd1984, 12'sd-1625}, {11'sd614, 12'sd-1338, 13'sd2544}},
{{9'sd210, 13'sd-2345, 13'sd2270}, {13'sd-2546, 11'sd597, 12'sd1178}, {12'sd1614, 13'sd2460, 13'sd-2161}},
{{9'sd231, 12'sd1684, 12'sd1111}, {11'sd940, 10'sd273, 11'sd-568}, {12'sd-1522, 12'sd-1849, 12'sd-1589}},
{{12'sd1392, 11'sd-627, 12'sd-1135}, {12'sd-1931, 11'sd-696, 12'sd-1097}, {12'sd-1401, 11'sd872, 10'sd-287}},
{{10'sd-320, 12'sd1570, 12'sd1280}, {11'sd1017, 10'sd-375, 12'sd1705}, {12'sd1031, 12'sd-1429, 12'sd1299}},
{{11'sd1003, 13'sd-3259, 13'sd-2550}, {11'sd-850, 8'sd-104, 12'sd1034}, {13'sd-2548, 6'sd-30, 11'sd623}},
{{13'sd2467, 11'sd-778, 11'sd722}, {12'sd-1929, 12'sd1936, 12'sd1739}, {12'sd1198, 12'sd-1159, 11'sd1017}},
{{11'sd795, 13'sd-2424, 11'sd733}, {10'sd-278, 5'sd14, 13'sd-2699}, {11'sd644, 13'sd-2417, 12'sd-1143}},
{{12'sd1379, 9'sd232, 12'sd1907}, {12'sd-1667, 11'sd816, 13'sd-2062}, {12'sd1244, 13'sd2142, 13'sd2084}},
{{11'sd929, 12'sd1526, 10'sd-388}, {12'sd1150, 11'sd-788, 11'sd-619}, {13'sd-2208, 11'sd-681, 13'sd-2797}},
{{10'sd-288, 13'sd2265, 12'sd1120}, {11'sd-992, 12'sd1618, 12'sd1940}, {13'sd2978, 13'sd2208, 10'sd375}}},
{
{{12'sd1170, 13'sd3041, 13'sd-2419}, {12'sd-2005, 12'sd1257, 10'sd279}, {10'sd275, 10'sd-399, 12'sd1126}},
{{13'sd2692, 5'sd11, 12'sd-1356}, {12'sd1738, 12'sd-1970, 9'sd217}, {13'sd2717, 12'sd-1121, 12'sd1925}},
{{13'sd-3533, 11'sd996, 11'sd-727}, {11'sd-779, 10'sd460, 11'sd-569}, {12'sd-1603, 12'sd-1599, 13'sd3188}},
{{9'sd-255, 13'sd2502, 12'sd1040}, {13'sd3003, 13'sd2929, 12'sd-1385}, {11'sd768, 9'sd233, 13'sd2639}},
{{10'sd-275, 12'sd1869, 12'sd1599}, {13'sd-2072, 13'sd2535, 10'sd269}, {10'sd-441, 9'sd-176, 9'sd207}},
{{12'sd1500, 11'sd533, 12'sd-1513}, {12'sd-1577, 13'sd2152, 12'sd1851}, {11'sd845, 12'sd1251, 12'sd1044}},
{{11'sd-836, 11'sd-977, 12'sd-2035}, {12'sd-1654, 12'sd1507, 11'sd535}, {12'sd-2026, 12'sd-1109, 11'sd882}},
{{13'sd-2183, 12'sd-1193, 7'sd-62}, {11'sd646, 11'sd-747, 10'sd273}, {12'sd1245, 13'sd2051, 11'sd997}},
{{11'sd-879, 11'sd944, 13'sd2327}, {13'sd-2212, 13'sd2963, 12'sd-1960}, {12'sd1292, 11'sd-901, 11'sd-785}},
{{12'sd1344, 12'sd-1118, 12'sd1265}, {13'sd-2780, 10'sd323, 12'sd-1621}, {13'sd2415, 10'sd-427, 7'sd32}},
{{14'sd4367, 13'sd2571, 13'sd-2247}, {10'sd-501, 11'sd589, 13'sd-2715}, {10'sd-421, 13'sd-2752, 12'sd-1948}},
{{13'sd-2205, 11'sd900, 12'sd1197}, {11'sd960, 11'sd859, 12'sd1420}, {13'sd2255, 12'sd1472, 13'sd2154}},
{{13'sd2550, 13'sd-2881, 13'sd2690}, {13'sd-3228, 8'sd125, 12'sd1106}, {13'sd-2097, 11'sd-926, 11'sd-536}},
{{13'sd2238, 10'sd471, 13'sd2097}, {11'sd-529, 11'sd-687, 12'sd-1783}, {10'sd-365, 13'sd-2219, 13'sd-2668}},
{{12'sd-1382, 10'sd-480, 10'sd-457}, {12'sd1349, 12'sd-1852, 13'sd-2345}, {10'sd462, 12'sd1271, 10'sd459}},
{{10'sd-430, 12'sd1471, 11'sd-623}, {11'sd1008, 12'sd-1193, 12'sd-1719}, {10'sd450, 6'sd22, 12'sd-1339}},
{{6'sd-24, 11'sd912, 12'sd1793}, {10'sd-309, 10'sd-268, 11'sd-771}, {13'sd2369, 11'sd-855, 3'sd-3}},
{{13'sd-3732, 12'sd-1353, 12'sd-1854}, {13'sd-2950, 11'sd668, 7'sd-59}, {13'sd3446, 12'sd1222, 11'sd-523}},
{{12'sd-1326, 13'sd-2535, 6'sd-31}, {13'sd-2215, 11'sd824, 10'sd-396}, {11'sd-836, 11'sd-538, 9'sd-182}},
{{12'sd-1159, 13'sd2500, 12'sd-1077}, {11'sd-921, 13'sd2479, 11'sd-646}, {10'sd345, 13'sd-2839, 12'sd-1034}},
{{10'sd362, 11'sd738, 9'sd-241}, {11'sd940, 11'sd-565, 13'sd-2473}, {10'sd-449, 13'sd2571, 13'sd2147}},
{{13'sd2219, 12'sd1879, 12'sd1771}, {11'sd-872, 12'sd1459, 10'sd409}, {13'sd2447, 13'sd-3237, 8'sd90}},
{{13'sd-2563, 12'sd-1521, 12'sd-1205}, {10'sd-257, 12'sd1184, 13'sd-2231}, {12'sd1532, 11'sd822, 8'sd108}},
{{13'sd2603, 13'sd-2444, 12'sd-1088}, {12'sd-1982, 11'sd649, 12'sd-1466}, {13'sd2108, 11'sd659, 12'sd-1568}},
{{11'sd718, 13'sd2362, 12'sd1102}, {12'sd-1551, 11'sd-581, 13'sd2373}, {10'sd352, 10'sd482, 13'sd3600}},
{{12'sd-1435, 11'sd-565, 10'sd-323}, {11'sd-549, 13'sd-2165, 11'sd-773}, {12'sd1682, 12'sd1084, 12'sd1525}},
{{13'sd2095, 12'sd-1172, 12'sd-1136}, {13'sd2119, 13'sd2805, 13'sd2551}, {12'sd1920, 11'sd596, 13'sd-2056}},
{{12'sd1411, 10'sd338, 11'sd779}, {12'sd1182, 12'sd1853, 12'sd-1030}, {12'sd-1152, 12'sd-1906, 13'sd2053}},
{{12'sd2018, 12'sd1523, 12'sd1196}, {12'sd-1879, 12'sd-1140, 12'sd-1204}, {12'sd1390, 11'sd-690, 11'sd1022}},
{{10'sd383, 12'sd-1721, 12'sd1971}, {12'sd-1427, 12'sd1121, 12'sd1285}, {12'sd-1449, 9'sd147, 12'sd1527}},
{{11'sd708, 13'sd-2288, 10'sd-361}, {13'sd2526, 11'sd-733, 13'sd2630}, {12'sd1939, 12'sd1624, 13'sd-2184}},
{{11'sd710, 13'sd-2308, 11'sd-887}, {9'sd248, 12'sd-1957, 12'sd-1115}, {11'sd-688, 13'sd2607, 10'sd437}},
{{13'sd2298, 13'sd-2237, 13'sd2193}, {12'sd-1605, 12'sd-1391, 10'sd-453}, {13'sd2210, 12'sd1212, 13'sd-2266}},
{{13'sd2786, 10'sd-433, 13'sd2745}, {12'sd-1532, 13'sd2176, 12'sd1878}, {12'sd-1186, 9'sd241, 13'sd-2164}},
{{12'sd1217, 13'sd2274, 11'sd794}, {13'sd-2423, 12'sd-1902, 11'sd-743}, {12'sd1446, 12'sd-1433, 13'sd-2380}},
{{12'sd-1652, 13'sd2370, 12'sd-1927}, {12'sd-1414, 13'sd2546, 9'sd-131}, {11'sd811, 13'sd2463, 12'sd1567}},
{{12'sd1966, 12'sd1902, 13'sd2367}, {13'sd3120, 12'sd-1477, 13'sd-2548}, {13'sd2110, 13'sd2957, 10'sd-328}},
{{12'sd-1770, 12'sd-1400, 13'sd-3122}, {12'sd-1819, 13'sd2906, 10'sd-511}, {9'sd-133, 13'sd2579, 13'sd-3206}},
{{12'sd1262, 12'sd1535, 12'sd-1712}, {12'sd-1745, 12'sd1360, 10'sd-458}, {12'sd-1314, 12'sd1159, 13'sd2096}},
{{12'sd-1405, 12'sd1271, 12'sd2042}, {13'sd-2171, 13'sd2292, 9'sd224}, {13'sd2798, 12'sd-1159, 12'sd1294}},
{{13'sd-2177, 12'sd-1659, 13'sd-2063}, {12'sd-1138, 10'sd340, 12'sd1893}, {12'sd1307, 11'sd705, 10'sd350}},
{{12'sd1105, 13'sd-2054, 11'sd-708}, {13'sd-2609, 11'sd898, 12'sd1042}, {4'sd7, 12'sd2032, 10'sd371}},
{{11'sd576, 12'sd-1469, 11'sd-677}, {10'sd392, 13'sd-2303, 13'sd-2281}, {12'sd1601, 12'sd1181, 11'sd662}},
{{11'sd-792, 13'sd-2053, 11'sd1009}, {12'sd-1772, 12'sd-2029, 12'sd1826}, {13'sd-3139, 10'sd316, 10'sd-347}},
{{11'sd654, 11'sd-562, 12'sd-2030}, {12'sd1661, 10'sd-438, 11'sd553}, {11'sd-621, 13'sd-2605, 13'sd-2308}},
{{11'sd-806, 10'sd498, 10'sd393}, {10'sd-482, 11'sd-611, 11'sd-822}, {12'sd-1868, 13'sd2300, 13'sd2564}},
{{13'sd-2300, 11'sd-954, 12'sd-1578}, {12'sd-2024, 11'sd571, 12'sd1241}, {12'sd2013, 12'sd-1237, 13'sd2504}},
{{12'sd1079, 12'sd1750, 11'sd711}, {11'sd594, 12'sd-1067, 11'sd732}, {11'sd-572, 12'sd-1393, 11'sd-838}},
{{12'sd2020, 12'sd1399, 12'sd-1506}, {13'sd2139, 12'sd-1594, 12'sd-1566}, {10'sd496, 12'sd-1877, 13'sd-2313}},
{{11'sd-650, 10'sd-504, 8'sd110}, {13'sd2603, 12'sd-1828, 12'sd-1646}, {11'sd725, 10'sd-339, 11'sd1023}},
{{13'sd-2599, 12'sd-1812, 11'sd-682}, {13'sd-2366, 10'sd-266, 13'sd2171}, {12'sd1380, 12'sd1066, 9'sd-138}},
{{11'sd981, 13'sd-2101, 11'sd830}, {12'sd1978, 13'sd-2300, 12'sd1244}, {12'sd-1590, 12'sd1433, 11'sd559}},
{{9'sd-165, 13'sd-2295, 11'sd515}, {7'sd-47, 12'sd-1518, 11'sd-744}, {13'sd3521, 8'sd93, 13'sd-2176}},
{{13'sd-2102, 13'sd-3020, 13'sd-2537}, {9'sd169, 13'sd-2472, 7'sd42}, {11'sd-692, 12'sd-1439, 13'sd-2726}},
{{13'sd-2450, 10'sd-480, 11'sd669}, {9'sd-246, 12'sd1068, 12'sd-1563}, {11'sd830, 13'sd-2570, 8'sd-101}},
{{12'sd-1218, 12'sd-1994, 12'sd-1236}, {12'sd-1117, 12'sd-1083, 12'sd-1559}, {12'sd-1643, 12'sd-1052, 8'sd110}},
{{11'sd1014, 12'sd1268, 11'sd-924}, {11'sd-697, 12'sd1109, 11'sd-917}, {12'sd-1606, 11'sd854, 12'sd1727}},
{{13'sd-3229, 12'sd-1860, 12'sd1142}, {12'sd-1357, 13'sd-2132, 10'sd346}, {12'sd1038, 12'sd1789, 13'sd2878}},
{{11'sd595, 12'sd-1913, 10'sd-256}, {12'sd1460, 9'sd173, 11'sd-949}, {10'sd355, 8'sd-76, 12'sd1409}},
{{13'sd-2457, 12'sd1836, 13'sd-2421}, {10'sd-389, 12'sd1053, 12'sd1325}, {11'sd-886, 12'sd1820, 12'sd1551}},
{{12'sd1270, 13'sd2814, 12'sd1342}, {13'sd-2504, 10'sd434, 13'sd-2388}, {13'sd-3016, 12'sd-1331, 11'sd-586}},
{{11'sd1005, 11'sd-1022, 11'sd-1013}, {11'sd-774, 10'sd-355, 5'sd-13}, {12'sd-1116, 11'sd671, 13'sd2073}},
{{11'sd763, 12'sd1273, 12'sd1424}, {10'sd-505, 13'sd-2659, 12'sd-1354}, {13'sd-2390, 11'sd621, 12'sd1352}},
{{9'sd-151, 9'sd158, 11'sd529}, {12'sd1433, 12'sd1939, 12'sd-2043}, {8'sd91, 11'sd-735, 12'sd1663}}},
{
{{12'sd-1051, 11'sd752, 8'sd125}, {8'sd68, 12'sd1687, 13'sd2618}, {13'sd-2361, 12'sd-1218, 12'sd1913}},
{{9'sd-152, 11'sd-1003, 7'sd-49}, {11'sd552, 13'sd3291, 11'sd863}, {13'sd-3522, 12'sd-1028, 13'sd3762}},
{{6'sd20, 12'sd1121, 12'sd1810}, {13'sd-2394, 12'sd1574, 12'sd-1726}, {13'sd-2488, 13'sd-2113, 13'sd-3559}},
{{12'sd-1625, 13'sd-2092, 12'sd1979}, {12'sd-2022, 12'sd-1575, 12'sd1368}, {12'sd-1222, 11'sd-647, 13'sd2372}},
{{13'sd-2151, 13'sd-2360, 12'sd-1229}, {12'sd1591, 10'sd387, 12'sd1247}, {12'sd1993, 13'sd-2205, 12'sd1407}},
{{12'sd-1068, 12'sd1222, 9'sd131}, {11'sd1023, 12'sd-1208, 12'sd1100}, {9'sd-148, 13'sd-2841, 12'sd-1675}},
{{13'sd-2364, 13'sd-3972, 9'sd250}, {13'sd-3359, 13'sd-4033, 13'sd-3402}, {12'sd1112, 12'sd1553, 12'sd1863}},
{{13'sd-3105, 13'sd-3053, 13'sd-3030}, {12'sd-1586, 12'sd1800, 12'sd-2021}, {11'sd-1007, 11'sd-630, 11'sd886}},
{{9'sd-239, 12'sd1841, 12'sd1368}, {12'sd-1260, 13'sd3553, 10'sd-325}, {10'sd-446, 12'sd1586, 6'sd-17}},
{{8'sd84, 11'sd-859, 12'sd-1496}, {12'sd-1075, 11'sd-910, 9'sd167}, {13'sd-2470, 12'sd-1285, 13'sd-2813}},
{{13'sd-3519, 6'sd-23, 12'sd-1857}, {14'sd-4949, 12'sd-1353, 6'sd-18}, {12'sd1416, 13'sd-3718, 11'sd905}},
{{11'sd941, 13'sd-2057, 12'sd-1539}, {13'sd2074, 7'sd-49, 13'sd2437}, {13'sd3275, 13'sd2863, 12'sd-1199}},
{{10'sd272, 13'sd-2293, 9'sd-246}, {12'sd-1414, 11'sd938, 12'sd1603}, {13'sd-2134, 6'sd31, 12'sd1850}},
{{13'sd-2634, 11'sd-788, 13'sd2174}, {12'sd1163, 12'sd-1871, 12'sd-1262}, {12'sd-1242, 9'sd-133, 10'sd488}},
{{13'sd-2540, 12'sd-1175, 11'sd-824}, {12'sd-1690, 13'sd-3495, 13'sd-2356}, {12'sd-1163, 13'sd-2214, 13'sd-2489}},
{{13'sd-2816, 13'sd-2259, 12'sd-1171}, {13'sd-3833, 13'sd-2666, 9'sd190}, {12'sd1306, 12'sd1085, 12'sd-1263}},
{{12'sd-1660, 13'sd-2109, 11'sd547}, {13'sd-3297, 11'sd911, 12'sd-1195}, {11'sd-602, 11'sd965, 13'sd2548}},
{{14'sd-6433, 13'sd-2434, 14'sd-4393}, {14'sd-4484, 12'sd-1596, 13'sd-4058}, {13'sd-3756, 12'sd-1464, 13'sd-2768}},
{{11'sd-871, 11'sd-717, 5'sd-8}, {12'sd1746, 12'sd-1347, 11'sd610}, {11'sd529, 10'sd-375, 11'sd-865}},
{{14'sd4457, 11'sd608, 10'sd393}, {13'sd3405, 12'sd1486, 8'sd-87}, {13'sd3075, 13'sd2939, 11'sd-994}},
{{13'sd3197, 11'sd982, 12'sd-1332}, {12'sd1784, 12'sd1911, 12'sd1925}, {12'sd-2036, 13'sd-2289, 12'sd-1634}},
{{11'sd747, 10'sd497, 12'sd1600}, {11'sd562, 13'sd-2653, 12'sd1570}, {13'sd-2095, 12'sd-1348, 11'sd520}},
{{12'sd-1548, 12'sd1567, 13'sd3144}, {13'sd-2974, 13'sd-2525, 12'sd1912}, {10'sd290, 13'sd-2160, 12'sd-1763}},
{{11'sd-1012, 12'sd-1245, 13'sd2604}, {12'sd-1319, 13'sd-2219, 12'sd-1094}, {13'sd-2586, 12'sd1246, 12'sd1236}},
{{9'sd243, 13'sd-2128, 11'sd-981}, {12'sd1900, 11'sd805, 9'sd-138}, {14'sd-4338, 13'sd-2664, 13'sd-3760}},
{{12'sd1194, 12'sd1877, 11'sd-817}, {13'sd2145, 12'sd-1419, 13'sd2221}, {10'sd-425, 13'sd2256, 13'sd2106}},
{{12'sd-1247, 12'sd1159, 12'sd-1795}, {8'sd65, 11'sd983, 12'sd1909}, {13'sd2072, 12'sd-1098, 12'sd-1318}},
{{12'sd-1328, 12'sd-1675, 9'sd181}, {12'sd-1923, 10'sd470, 9'sd224}, {12'sd1902, 11'sd-604, 11'sd-750}},
{{10'sd-412, 13'sd-2991, 12'sd-1862}, {13'sd-2967, 13'sd-2079, 9'sd248}, {13'sd2668, 12'sd-1734, 13'sd-2269}},
{{12'sd-1164, 13'sd-2826, 11'sd-902}, {11'sd-831, 12'sd1899, 11'sd-660}, {13'sd2448, 12'sd1128, 9'sd-219}},
{{11'sd546, 11'sd-779, 11'sd814}, {10'sd-333, 13'sd-2172, 12'sd-1626}, {12'sd-1336, 9'sd-242, 13'sd2144}},
{{11'sd981, 13'sd2155, 12'sd1092}, {13'sd-2329, 10'sd-449, 10'sd-322}, {12'sd-1751, 12'sd-1494, 13'sd2716}},
{{13'sd2824, 11'sd-1006, 10'sd-359}, {12'sd-1352, 13'sd2476, 11'sd-533}, {13'sd-2767, 10'sd-273, 13'sd2632}},
{{13'sd4032, 10'sd-489, 13'sd2846}, {10'sd-343, 12'sd-1816, 11'sd884}, {12'sd1307, 12'sd1460, 13'sd-2570}},
{{12'sd1437, 13'sd-2857, 12'sd1691}, {11'sd-801, 11'sd-637, 11'sd-773}, {13'sd3422, 13'sd2373, 11'sd577}},
{{12'sd-1229, 12'sd1156, 11'sd886}, {10'sd-410, 12'sd-1526, 11'sd-630}, {13'sd3109, 12'sd1294, 12'sd1144}},
{{13'sd3012, 13'sd2978, 13'sd2615}, {12'sd1716, 12'sd-1366, 13'sd3578}, {12'sd1963, 10'sd-416, 11'sd-596}},
{{13'sd-2749, 13'sd-3890, 10'sd-283}, {14'sd-4328, 11'sd-721, 13'sd3459}, {11'sd-620, 12'sd-1414, 13'sd3619}},
{{12'sd-1202, 10'sd-262, 13'sd-2117}, {12'sd-1987, 11'sd949, 7'sd-34}, {12'sd-1625, 13'sd2123, 12'sd-1739}},
{{8'sd120, 13'sd-2648, 10'sd-257}, {5'sd-15, 10'sd445, 13'sd-2095}, {12'sd1102, 12'sd-1070, 12'sd1889}},
{{13'sd-3348, 13'sd-2415, 11'sd-732}, {13'sd-3553, 13'sd-2105, 13'sd2256}, {13'sd-3472, 10'sd-264, 13'sd2123}},
{{10'sd-399, 12'sd-1688, 12'sd-1735}, {11'sd880, 12'sd1756, 13'sd2188}, {13'sd-2376, 11'sd-572, 13'sd2564}},
{{11'sd-854, 12'sd1180, 13'sd2236}, {12'sd-1605, 11'sd624, 11'sd569}, {13'sd2935, 10'sd-483, 6'sd-27}},
{{12'sd2034, 12'sd1253, 11'sd783}, {13'sd2453, 13'sd3273, 9'sd-167}, {11'sd732, 10'sd-272, 10'sd-290}},
{{13'sd2101, 8'sd72, 13'sd-2445}, {13'sd-2750, 8'sd-124, 13'sd-2621}, {11'sd-939, 11'sd-712, 11'sd-724}},
{{7'sd49, 13'sd2834, 8'sd-84}, {10'sd396, 12'sd1156, 11'sd-993}, {12'sd1164, 13'sd-3963, 14'sd-4138}},
{{14'sd-4560, 11'sd-1018, 9'sd-139}, {14'sd-4769, 11'sd989, 13'sd-3146}, {13'sd-2375, 12'sd-1608, 13'sd-2259}},
{{12'sd-1884, 10'sd379, 12'sd1822}, {10'sd-326, 6'sd-20, 11'sd749}, {12'sd-1235, 8'sd-70, 3'sd2}},
{{11'sd-959, 12'sd1129, 12'sd-1339}, {11'sd-810, 12'sd-1426, 12'sd1338}, {13'sd2282, 10'sd-496, 8'sd74}},
{{13'sd-2594, 8'sd64, 11'sd1003}, {7'sd42, 13'sd-2072, 12'sd-1819}, {12'sd1768, 11'sd-656, 10'sd411}},
{{11'sd-803, 12'sd1325, 13'sd-2546}, {9'sd-158, 11'sd939, 11'sd-742}, {12'sd-1548, 11'sd573, 12'sd-1066}},
{{13'sd2305, 13'sd2093, 10'sd-416}, {11'sd659, 12'sd1085, 12'sd1417}, {8'sd-89, 11'sd904, 12'sd1369}},
{{11'sd-862, 14'sd-4453, 12'sd1622}, {12'sd-1801, 9'sd226, 11'sd707}, {13'sd-3723, 12'sd-1734, 12'sd-2000}},
{{11'sd987, 13'sd2166, 13'sd3089}, {12'sd-1118, 12'sd1652, 9'sd-183}, {11'sd884, 12'sd1140, 12'sd1864}},
{{11'sd-634, 11'sd735, 13'sd2780}, {10'sd380, 12'sd1300, 13'sd-2456}, {13'sd-2387, 12'sd-1609, 12'sd1602}},
{{13'sd2545, 12'sd-1271, 13'sd3007}, {12'sd-1478, 13'sd-2481, 13'sd2332}, {12'sd1601, 10'sd281, 12'sd-1499}},
{{11'sd997, 12'sd1158, 13'sd2491}, {12'sd-1250, 13'sd-2985, 12'sd1438}, {12'sd-1660, 13'sd-3136, 12'sd1799}},
{{12'sd-1109, 12'sd1437, 12'sd-1048}, {10'sd294, 10'sd-299, 11'sd736}, {13'sd-2890, 10'sd-358, 11'sd940}},
{{12'sd1841, 9'sd236, 12'sd-1845}, {8'sd-122, 13'sd2588, 12'sd-1050}, {13'sd-3725, 13'sd-3104, 12'sd-1982}},
{{12'sd-1546, 11'sd-576, 13'sd-3040}, {11'sd-808, 9'sd-236, 13'sd-2605}, {13'sd2220, 12'sd1902, 13'sd-2159}},
{{11'sd704, 9'sd-202, 11'sd-574}, {13'sd3859, 10'sd-275, 13'sd2595}, {13'sd2553, 13'sd2100, 11'sd-885}},
{{12'sd-1711, 11'sd-977, 13'sd-2939}, {12'sd1126, 12'sd1131, 12'sd-1923}, {13'sd2384, 12'sd1506, 13'sd2328}},
{{8'sd-69, 14'sd4306, 11'sd676}, {12'sd1900, 14'sd4275, 13'sd2738}, {12'sd1111, 13'sd2247, 11'sd857}},
{{7'sd37, 12'sd1958, 12'sd-1483}, {13'sd3082, 10'sd-426, 10'sd408}, {11'sd-981, 5'sd10, 12'sd-1061}}},
{
{{14'sd4631, 13'sd2279, 12'sd-1715}, {13'sd2279, 12'sd1871, 13'sd-3193}, {11'sd-805, 11'sd833, 11'sd-764}},
{{11'sd-782, 13'sd2684, 13'sd2369}, {11'sd-946, 13'sd-2726, 13'sd-2102}, {13'sd2281, 12'sd-1100, 13'sd-2814}},
{{13'sd-2171, 13'sd2931, 11'sd-906}, {12'sd-1744, 10'sd445, 10'sd263}, {13'sd-3093, 12'sd-1522, 10'sd386}},
{{8'sd-123, 13'sd-3014, 13'sd2460}, {13'sd2382, 9'sd132, 10'sd388}, {11'sd-914, 11'sd-729, 12'sd1299}},
{{13'sd3341, 12'sd-1187, 13'sd2850}, {11'sd518, 12'sd1230, 13'sd2810}, {13'sd2207, 12'sd1617, 13'sd2176}},
{{13'sd2076, 11'sd-768, 9'sd-233}, {12'sd1908, 11'sd-581, 13'sd2337}, {12'sd-1113, 10'sd-508, 10'sd477}},
{{11'sd850, 12'sd-1376, 12'sd-1857}, {11'sd725, 6'sd28, 13'sd-2560}, {13'sd2655, 11'sd-758, 8'sd127}},
{{10'sd-274, 11'sd-793, 12'sd-1053}, {13'sd2062, 13'sd-2982, 12'sd-1274}, {10'sd-311, 12'sd1024, 10'sd-393}},
{{11'sd-714, 13'sd2567, 13'sd2301}, {12'sd1153, 12'sd-1122, 11'sd-923}, {12'sd-1958, 11'sd-898, 12'sd1040}},
{{11'sd789, 12'sd2029, 12'sd1140}, {12'sd-1641, 12'sd-1254, 11'sd765}, {12'sd1869, 13'sd-2809, 13'sd-2982}},
{{13'sd-3206, 11'sd553, 11'sd-730}, {12'sd-1765, 13'sd-2830, 11'sd919}, {14'sd4800, 13'sd2286, 14'sd5388}},
{{9'sd-178, 12'sd1130, 11'sd759}, {12'sd-1272, 13'sd-2219, 12'sd-1074}, {9'sd206, 11'sd-549, 12'sd-1436}},
{{12'sd-1418, 13'sd2801, 13'sd-3712}, {12'sd1117, 13'sd2975, 11'sd-539}, {12'sd-1878, 13'sd2583, 9'sd228}},
{{10'sd-402, 13'sd-2310, 10'sd344}, {12'sd-1411, 13'sd2347, 11'sd-972}, {10'sd463, 12'sd-1819, 12'sd1609}},
{{12'sd1318, 13'sd2061, 11'sd549}, {11'sd976, 12'sd1133, 13'sd2778}, {11'sd-827, 12'sd-1540, 13'sd2486}},
{{12'sd1975, 11'sd-724, 9'sd222}, {12'sd1343, 11'sd-764, 12'sd1117}, {13'sd3121, 11'sd-763, 13'sd2717}},
{{12'sd1443, 10'sd-356, 12'sd1754}, {12'sd-1995, 13'sd3410, 12'sd1979}, {11'sd871, 13'sd3729, 10'sd441}},
{{10'sd-304, 12'sd1710, 10'sd-299}, {13'sd2395, 12'sd1336, 12'sd1994}, {13'sd3802, 13'sd3576, 10'sd-304}},
{{12'sd-1373, 11'sd656, 11'sd-934}, {13'sd2939, 12'sd-2043, 10'sd370}, {12'sd-1159, 8'sd-90, 13'sd-2323}},
{{7'sd-41, 12'sd-1305, 12'sd-1184}, {2'sd1, 10'sd-298, 9'sd201}, {12'sd-1639, 12'sd1867, 13'sd-2590}},
{{7'sd53, 13'sd2487, 11'sd-939}, {12'sd-1519, 10'sd-370, 12'sd1179}, {9'sd-155, 12'sd1460, 12'sd1081}},
{{12'sd-1765, 13'sd-2945, 10'sd-432}, {13'sd-2975, 9'sd-172, 8'sd118}, {10'sd-275, 8'sd-77, 10'sd338}},
{{11'sd610, 8'sd91, 10'sd292}, {12'sd1617, 12'sd-1964, 11'sd-526}, {12'sd1813, 13'sd-2342, 10'sd-279}},
{{12'sd-1964, 11'sd842, 13'sd2343}, {11'sd649, 13'sd-2990, 12'sd1465}, {11'sd904, 13'sd-2139, 12'sd1557}},
{{14'sd4502, 14'sd4573, 12'sd1085}, {11'sd-519, 14'sd4247, 13'sd-2204}, {11'sd637, 13'sd-2779, 13'sd-3242}},
{{13'sd2350, 12'sd-1158, 12'sd1518}, {12'sd1127, 10'sd-348, 10'sd-454}, {3'sd3, 13'sd2370, 13'sd-2082}},
{{12'sd1052, 12'sd-1142, 12'sd-1678}, {12'sd-1244, 12'sd-1759, 12'sd1038}, {10'sd464, 10'sd351, 11'sd974}},
{{8'sd70, 13'sd-2303, 13'sd2509}, {12'sd1698, 12'sd1756, 12'sd1762}, {13'sd2623, 13'sd-2333, 11'sd961}},
{{12'sd-1091, 11'sd-542, 13'sd-2068}, {9'sd149, 13'sd2344, 13'sd-2052}, {13'sd2420, 11'sd-969, 13'sd3249}},
{{8'sd-74, 13'sd-3521, 13'sd-2140}, {11'sd1022, 12'sd-1742, 13'sd3066}, {9'sd-129, 12'sd1831, 10'sd-470}},
{{10'sd433, 12'sd1282, 12'sd1769}, {10'sd318, 13'sd2691, 12'sd1055}, {13'sd-2465, 12'sd-1443, 11'sd-541}},
{{13'sd2880, 9'sd139, 11'sd571}, {12'sd-1956, 12'sd-1603, 13'sd-2319}, {12'sd-1722, 12'sd1962, 12'sd-1864}},
{{11'sd965, 12'sd-1811, 12'sd-1562}, {10'sd363, 12'sd1399, 13'sd-2845}, {13'sd2280, 11'sd809, 10'sd-477}},
{{13'sd-2549, 11'sd884, 13'sd2260}, {10'sd-480, 11'sd912, 12'sd1499}, {10'sd409, 12'sd-1222, 10'sd386}},
{{12'sd-1269, 12'sd1459, 10'sd305}, {9'sd218, 12'sd1232, 9'sd139}, {11'sd918, 12'sd1981, 7'sd-44}},
{{13'sd2402, 13'sd-2431, 13'sd2238}, {11'sd593, 12'sd1923, 12'sd-1365}, {12'sd-1080, 12'sd1895, 12'sd-1539}},
{{10'sd496, 12'sd1893, 13'sd3691}, {12'sd2022, 11'sd810, 12'sd1663}, {13'sd-2141, 13'sd2239, 10'sd-428}},
{{13'sd3324, 11'sd-538, 13'sd2292}, {12'sd1247, 13'sd2606, 11'sd-735}, {13'sd4020, 11'sd-678, 12'sd1841}},
{{12'sd1441, 12'sd1252, 12'sd1673}, {10'sd280, 13'sd-2136, 10'sd-451}, {13'sd3477, 11'sd570, 10'sd350}},
{{12'sd1330, 11'sd908, 14'sd-4109}, {9'sd233, 11'sd1005, 8'sd98}, {13'sd2312, 11'sd738, 9'sd219}},
{{7'sd63, 13'sd3116, 12'sd-1443}, {13'sd-2501, 13'sd3334, 13'sd-2857}, {11'sd-823, 9'sd159, 10'sd-319}},
{{12'sd1164, 9'sd216, 7'sd59}, {12'sd1861, 10'sd319, 4'sd-6}, {8'sd81, 10'sd444, 11'sd-997}},
{{12'sd-1233, 13'sd-3797, 13'sd-3045}, {13'sd2538, 12'sd1518, 12'sd1117}, {11'sd-701, 12'sd-1141, 10'sd-507}},
{{10'sd362, 9'sd152, 13'sd-2337}, {13'sd-2804, 12'sd-1742, 13'sd-2082}, {14'sd-4252, 13'sd-3923, 12'sd-1098}},
{{13'sd-2477, 9'sd-132, 12'sd-1466}, {11'sd939, 12'sd1514, 12'sd1844}, {12'sd-1709, 12'sd1495, 10'sd-336}},
{{12'sd-1281, 13'sd2951, 12'sd1849}, {13'sd-2646, 11'sd-970, 12'sd-1101}, {12'sd-1670, 10'sd403, 8'sd85}},
{{12'sd1887, 10'sd278, 12'sd-1433}, {9'sd-138, 12'sd-1079, 7'sd-60}, {12'sd-1693, 12'sd1322, 12'sd1097}},
{{12'sd-1850, 12'sd2045, 12'sd-1326}, {10'sd256, 9'sd240, 11'sd-750}, {11'sd-959, 12'sd1369, 10'sd277}},
{{8'sd-66, 12'sd1198, 9'sd238}, {11'sd-804, 6'sd-19, 8'sd117}, {13'sd-2847, 12'sd1305, 12'sd-1841}},
{{12'sd1991, 12'sd-1481, 12'sd-1354}, {11'sd539, 13'sd2321, 12'sd1925}, {9'sd141, 12'sd1893, 9'sd-153}},
{{9'sd155, 12'sd-1888, 11'sd901}, {12'sd-1098, 12'sd1425, 12'sd-1275}, {9'sd-196, 10'sd-507, 9'sd-230}},
{{13'sd2549, 11'sd797, 13'sd-2207}, {12'sd-1257, 11'sd-987, 10'sd-303}, {13'sd2372, 10'sd-263, 13'sd2520}},
{{10'sd-339, 10'sd328, 13'sd2896}, {12'sd-1527, 12'sd1204, 11'sd908}, {11'sd581, 13'sd3162, 14'sd6031}},
{{13'sd2422, 12'sd-1956, 12'sd-2034}, {11'sd718, 13'sd2522, 13'sd-2661}, {11'sd-726, 12'sd1607, 7'sd45}},
{{12'sd-1374, 11'sd789, 13'sd-2250}, {12'sd1406, 12'sd-1119, 12'sd-1236}, {12'sd1504, 13'sd-2377, 9'sd174}},
{{12'sd1640, 11'sd-848, 11'sd-1008}, {12'sd-1123, 13'sd2508, 12'sd-1498}, {12'sd-1566, 9'sd-221, 11'sd-636}},
{{11'sd-618, 12'sd1097, 12'sd-1898}, {13'sd-2889, 12'sd-1731, 7'sd-60}, {13'sd-2754, 12'sd1852, 13'sd2711}},
{{10'sd472, 8'sd110, 12'sd-1188}, {13'sd2102, 12'sd-1047, 11'sd-646}, {8'sd-78, 12'sd-1085, 13'sd-2203}},
{{13'sd2454, 12'sd1417, 13'sd-2167}, {11'sd850, 12'sd-1704, 11'sd1023}, {13'sd2105, 9'sd-250, 13'sd-2811}},
{{13'sd-2588, 13'sd-2766, 12'sd1332}, {13'sd-2113, 12'sd1660, 11'sd-740}, {8'sd-82, 12'sd1420, 12'sd1477}},
{{13'sd-2180, 13'sd-2431, 13'sd2312}, {13'sd2895, 7'sd48, 13'sd-3731}, {13'sd-2082, 10'sd-487, 13'sd-2637}},
{{12'sd-1228, 12'sd-1115, 11'sd-849}, {10'sd378, 12'sd-1786, 12'sd1487}, {10'sd269, 10'sd410, 12'sd-1352}},
{{12'sd1089, 10'sd-441, 12'sd-1157}, {9'sd-200, 11'sd-985, 12'sd1528}, {13'sd-2681, 13'sd2209, 11'sd-889}},
{{13'sd2526, 12'sd1582, 13'sd-2405}, {12'sd-1723, 12'sd-1754, 12'sd-1921}, {13'sd2323, 12'sd1863, 13'sd-3467}}},
{
{{12'sd1803, 9'sd140, 12'sd-1076}, {13'sd-2441, 10'sd338, 13'sd-2767}, {11'sd593, 12'sd1227, 13'sd-2563}},
{{13'sd2345, 12'sd2003, 12'sd-1509}, {13'sd2520, 12'sd2028, 12'sd1711}, {9'sd253, 11'sd-544, 13'sd2546}},
{{13'sd2284, 10'sd475, 14'sd4785}, {13'sd3029, 12'sd1833, 12'sd1985}, {13'sd2164, 9'sd151, 12'sd-1469}},
{{12'sd1079, 10'sd397, 11'sd-688}, {10'sd400, 12'sd-1333, 13'sd-3694}, {11'sd-1006, 13'sd-2500, 9'sd190}},
{{13'sd3734, 11'sd-878, 12'sd-1706}, {13'sd3013, 10'sd-499, 11'sd737}, {12'sd1212, 14'sd-4241, 13'sd-2894}},
{{13'sd-2559, 12'sd-1035, 13'sd-2858}, {6'sd28, 13'sd-2504, 6'sd-18}, {7'sd49, 11'sd978, 11'sd800}},
{{12'sd-1294, 11'sd633, 11'sd-711}, {13'sd2253, 13'sd2724, 10'sd430}, {10'sd354, 13'sd2184, 12'sd-1457}},
{{7'sd62, 12'sd1133, 12'sd1311}, {12'sd1832, 12'sd-2043, 12'sd-1342}, {10'sd-288, 13'sd-2453, 10'sd349}},
{{12'sd1751, 13'sd-2254, 11'sd633}, {10'sd464, 12'sd1533, 12'sd-1837}, {11'sd895, 12'sd1986, 12'sd-2035}},
{{12'sd1195, 11'sd619, 14'sd-4635}, {13'sd3887, 13'sd2525, 11'sd-595}, {12'sd1563, 10'sd488, 13'sd2080}},
{{14'sd-5735, 10'sd-341, 13'sd2224}, {13'sd-3351, 12'sd-1895, 13'sd3138}, {13'sd-3129, 13'sd-2954, 10'sd-511}},
{{12'sd1877, 12'sd-1153, 12'sd1028}, {12'sd-1605, 12'sd1903, 11'sd515}, {12'sd1112, 11'sd999, 5'sd14}},
{{12'sd1817, 14'sd6079, 13'sd2215}, {13'sd3724, 13'sd3959, 11'sd-664}, {11'sd960, 10'sd478, 13'sd3838}},
{{13'sd2500, 11'sd-977, 5'sd-9}, {12'sd-1593, 13'sd-2782, 13'sd-3197}, {12'sd-1268, 12'sd1436, 12'sd-1580}},
{{13'sd-2422, 10'sd455, 13'sd2497}, {13'sd-2455, 13'sd2167, 11'sd-633}, {12'sd1197, 13'sd-2931, 9'sd-254}},
{{12'sd1271, 12'sd1070, 11'sd-646}, {13'sd2080, 10'sd-411, 12'sd-1842}, {10'sd-404, 12'sd1065, 11'sd-520}},
{{13'sd2598, 11'sd-895, 13'sd-2576}, {10'sd319, 11'sd619, 12'sd1285}, {12'sd1796, 13'sd2374, 11'sd-719}},
{{14'sd6244, 11'sd753, 13'sd-2861}, {14'sd4115, 13'sd3239, 11'sd-832}, {10'sd400, 13'sd-2132, 11'sd-850}},
{{6'sd18, 11'sd758, 13'sd-2938}, {6'sd-25, 10'sd329, 12'sd1856}, {10'sd-342, 12'sd-1279, 13'sd-2760}},
{{12'sd1068, 13'sd-3042, 12'sd-1441}, {12'sd1448, 12'sd-1792, 12'sd1123}, {3'sd3, 14'sd-4525, 9'sd-230}},
{{10'sd504, 13'sd-2938, 12'sd1289}, {13'sd2269, 12'sd1053, 12'sd-1223}, {11'sd-568, 10'sd506, 13'sd2578}},
{{12'sd1350, 13'sd2734, 12'sd1893}, {12'sd-1278, 12'sd1344, 11'sd-651}, {11'sd-1010, 13'sd-2091, 12'sd-1142}},
{{12'sd-1030, 13'sd-3254, 11'sd839}, {12'sd-1979, 13'sd-2488, 11'sd-819}, {13'sd-2118, 11'sd872, 12'sd1510}},
{{11'sd-701, 12'sd1961, 12'sd-1106}, {9'sd190, 7'sd54, 12'sd-1295}, {12'sd-1096, 10'sd494, 13'sd2135}},
{{10'sd-352, 12'sd-1270, 10'sd-307}, {11'sd-786, 13'sd-2523, 13'sd-2207}, {14'sd4147, 11'sd551, 13'sd3993}},
{{9'sd-150, 12'sd1768, 13'sd2539}, {12'sd1076, 12'sd-1237, 11'sd822}, {11'sd-846, 10'sd272, 13'sd-3040}},
{{13'sd3010, 13'sd2197, 10'sd-292}, {12'sd-1303, 4'sd5, 13'sd-3517}, {12'sd-1232, 13'sd-2149, 12'sd-1474}},
{{13'sd2435, 11'sd552, 13'sd-2592}, {10'sd466, 10'sd-402, 13'sd-3796}, {13'sd2815, 12'sd-1560, 11'sd-956}},
{{13'sd2241, 12'sd1810, 12'sd1252}, {7'sd52, 11'sd654, 13'sd3743}, {12'sd-1450, 11'sd849, 13'sd2935}},
{{13'sd3720, 12'sd-1105, 10'sd268}, {13'sd2795, 12'sd1565, 12'sd1961}, {12'sd-1203, 12'sd-1794, 12'sd1885}},
{{12'sd-1857, 13'sd-3323, 13'sd2257}, {13'sd-2105, 12'sd1220, 13'sd3306}, {12'sd-1678, 11'sd984, 10'sd395}},
{{13'sd-3229, 10'sd-460, 13'sd-3053}, {12'sd-1969, 8'sd88, 11'sd648}, {11'sd748, 13'sd-2845, 9'sd-247}},
{{12'sd1309, 11'sd-815, 11'sd700}, {12'sd1814, 13'sd2668, 11'sd-908}, {9'sd242, 11'sd-691, 14'sd4224}},
{{12'sd-1579, 13'sd-3156, 13'sd-4083}, {12'sd-1314, 12'sd-1899, 12'sd-1566}, {13'sd-3192, 12'sd1363, 13'sd2415}},
{{10'sd-281, 13'sd3231, 12'sd1255}, {13'sd-2322, 11'sd-755, 9'sd180}, {11'sd901, 8'sd113, 11'sd-597}},
{{11'sd587, 11'sd639, 12'sd-1160}, {8'sd-99, 11'sd-563, 11'sd654}, {13'sd2720, 12'sd-1601, 11'sd-966}},
{{12'sd1870, 10'sd-390, 10'sd347}, {10'sd-397, 12'sd1062, 9'sd202}, {11'sd-908, 13'sd2487, 12'sd-1547}},
{{14'sd4689, 12'sd-1702, 11'sd987}, {13'sd3767, 10'sd292, 12'sd-1168}, {12'sd-1691, 13'sd-3931, 13'sd-3061}},
{{13'sd-2211, 6'sd29, 13'sd2848}, {12'sd1221, 12'sd-1156, 11'sd-876}, {10'sd428, 10'sd-293, 12'sd-1430}},
{{12'sd1049, 10'sd374, 14'sd4319}, {8'sd-98, 13'sd3352, 9'sd162}, {13'sd-2357, 12'sd-1638, 13'sd-2742}},
{{11'sd-552, 12'sd-1442, 13'sd2079}, {12'sd1436, 12'sd-1036, 8'sd64}, {12'sd-1313, 12'sd1097, 10'sd-339}},
{{12'sd1804, 1'sd0, 12'sd1506}, {12'sd1534, 13'sd2256, 11'sd750}, {10'sd-293, 11'sd803, 10'sd343}},
{{13'sd-2188, 12'sd1648, 12'sd1267}, {13'sd-3259, 13'sd-2361, 11'sd-734}, {12'sd-1340, 13'sd-2595, 13'sd-3668}},
{{13'sd-2209, 12'sd1283, 13'sd2690}, {12'sd1090, 13'sd-2977, 11'sd614}, {13'sd-3229, 11'sd-787, 12'sd-1884}},
{{12'sd1200, 5'sd-11, 11'sd888}, {13'sd-2056, 12'sd1740, 11'sd-712}, {7'sd56, 11'sd806, 13'sd2574}},
{{10'sd-463, 13'sd-2639, 12'sd-1577}, {12'sd1048, 11'sd684, 13'sd2112}, {9'sd223, 13'sd2694, 12'sd1848}},
{{10'sd378, 11'sd-800, 12'sd-1870}, {14'sd4136, 12'sd1944, 13'sd2464}, {11'sd-829, 11'sd728, 13'sd3172}},
{{9'sd-213, 4'sd-6, 12'sd-1121}, {13'sd-2211, 9'sd-188, 12'sd1591}, {11'sd682, 8'sd86, 10'sd452}},
{{11'sd1018, 13'sd3350, 12'sd-1339}, {10'sd-344, 13'sd-2993, 13'sd-3354}, {12'sd1141, 11'sd531, 13'sd-2549}},
{{13'sd2393, 13'sd4040, 13'sd2470}, {11'sd-875, 12'sd1358, 12'sd-1037}, {12'sd1167, 13'sd2118, 13'sd3218}},
{{12'sd1452, 13'sd3986, 13'sd2978}, {12'sd-1158, 10'sd299, 13'sd-3313}, {12'sd-1405, 12'sd-1612, 10'sd-479}},
{{9'sd-164, 12'sd-1518, 13'sd-2673}, {12'sd-1463, 12'sd-1316, 11'sd800}, {13'sd-2094, 12'sd1720, 13'sd2562}},
{{10'sd-311, 13'sd-2061, 13'sd2882}, {12'sd-1076, 13'sd2650, 13'sd-2132}, {13'sd-2493, 11'sd800, 10'sd402}},
{{10'sd398, 12'sd-1382, 11'sd993}, {11'sd-655, 10'sd423, 13'sd3214}, {9'sd209, 11'sd-543, 13'sd2157}},
{{11'sd-996, 13'sd-2225, 12'sd-1809}, {13'sd-2235, 8'sd-74, 10'sd384}, {12'sd1385, 13'sd-2399, 12'sd1636}},
{{13'sd-2943, 13'sd-2191, 12'sd-1292}, {10'sd-357, 12'sd-1472, 10'sd-325}, {7'sd50, 13'sd2858, 13'sd2522}},
{{11'sd-882, 12'sd-1254, 11'sd-1023}, {12'sd1119, 12'sd1505, 9'sd220}, {12'sd1745, 12'sd2032, 14'sd4674}},
{{11'sd-764, 12'sd1630, 12'sd-1050}, {13'sd2089, 12'sd-1583, 10'sd376}, {12'sd1245, 12'sd1122, 11'sd-635}},
{{11'sd-967, 12'sd-1995, 10'sd-440}, {13'sd-3894, 11'sd-801, 11'sd-1012}, {13'sd-3821, 13'sd-2896, 13'sd-2390}},
{{10'sd-319, 8'sd-84, 12'sd-1741}, {11'sd693, 12'sd1557, 11'sd825}, {10'sd-421, 13'sd2052, 13'sd-2493}},
{{10'sd-300, 12'sd1449, 11'sd-607}, {11'sd523, 12'sd1923, 13'sd-2552}, {12'sd1290, 10'sd499, 13'sd-3030}},
{{13'sd3332, 13'sd2859, 11'sd576}, {13'sd2227, 12'sd1780, 12'sd1738}, {13'sd2210, 9'sd-171, 12'sd1704}},
{{11'sd800, 7'sd53, 12'sd-1203}, {12'sd1437, 14'sd-4824, 12'sd-1147}, {11'sd587, 11'sd591, 10'sd-385}},
{{12'sd1466, 11'sd802, 12'sd1717}, {12'sd-1262, 12'sd-1393, 11'sd590}, {12'sd-1695, 11'sd699, 13'sd-3465}}},
{
{{10'sd298, 12'sd-1542, 13'sd3134}, {13'sd-2322, 12'sd1500, 13'sd4028}, {12'sd1398, 12'sd1077, 8'sd75}},
{{12'sd1172, 13'sd-2066, 13'sd-3989}, {12'sd-1759, 12'sd1224, 11'sd-1009}, {11'sd839, 13'sd3844, 13'sd-2307}},
{{11'sd-547, 11'sd569, 10'sd261}, {13'sd-2384, 13'sd-2543, 12'sd1459}, {9'sd-150, 11'sd-601, 13'sd2510}},
{{10'sd-466, 13'sd2456, 12'sd-1730}, {12'sd-1414, 11'sd-971, 13'sd2132}, {8'sd100, 11'sd942, 13'sd2449}},
{{13'sd-3174, 12'sd1162, 11'sd909}, {12'sd-1821, 13'sd2408, 9'sd198}, {12'sd1142, 13'sd2517, 12'sd1729}},
{{12'sd-1816, 10'sd-389, 13'sd-3466}, {13'sd2938, 9'sd-170, 13'sd-3102}, {12'sd1747, 11'sd646, 12'sd-1942}},
{{11'sd-647, 11'sd-666, 11'sd604}, {12'sd-1566, 13'sd-2699, 13'sd-2332}, {9'sd246, 8'sd-79, 11'sd1005}},
{{13'sd-2284, 13'sd-2130, 11'sd640}, {8'sd109, 12'sd-2016, 13'sd2484}, {12'sd-2029, 12'sd1742, 12'sd-1095}},
{{11'sd772, 8'sd-104, 12'sd-1781}, {13'sd3235, 13'sd2850, 11'sd1019}, {12'sd1458, 12'sd-1947, 11'sd577}},
{{11'sd929, 12'sd1662, 13'sd-3647}, {11'sd-634, 10'sd381, 13'sd-2771}, {13'sd-3860, 12'sd1542, 10'sd281}},
{{13'sd-3905, 11'sd-638, 14'sd4880}, {11'sd855, 10'sd400, 12'sd1685}, {13'sd-3108, 8'sd-104, 13'sd3260}},
{{7'sd48, 11'sd534, 11'sd-521}, {10'sd299, 12'sd-1490, 12'sd-1112}, {13'sd-2112, 13'sd2897, 12'sd1403}},
{{13'sd3151, 9'sd223, 8'sd-65}, {13'sd2147, 13'sd2224, 12'sd-1604}, {14'sd5057, 11'sd-530, 11'sd655}},
{{8'sd-122, 9'sd-200, 13'sd-2175}, {10'sd-442, 12'sd-1939, 11'sd-931}, {12'sd1437, 9'sd-238, 11'sd597}},
{{13'sd-2471, 13'sd-2609, 6'sd-26}, {7'sd36, 12'sd2044, 12'sd-1656}, {7'sd43, 12'sd-1753, 11'sd916}},
{{11'sd546, 13'sd-2121, 12'sd-1741}, {12'sd1042, 11'sd-786, 12'sd-1741}, {12'sd1795, 13'sd2295, 10'sd440}},
{{9'sd200, 12'sd1299, 13'sd-3028}, {13'sd2358, 13'sd2538, 10'sd451}, {12'sd-1442, 9'sd-147, 13'sd3100}},
{{13'sd-3327, 12'sd-1089, 14'sd-6652}, {11'sd883, 13'sd-2354, 11'sd552}, {12'sd-1498, 10'sd470, 13'sd-2929}},
{{12'sd1939, 11'sd-610, 13'sd2626}, {11'sd-771, 12'sd1451, 11'sd1003}, {13'sd-2138, 11'sd-898, 12'sd1152}},
{{12'sd-1369, 10'sd294, 14'sd-5217}, {9'sd-185, 12'sd1306, 13'sd-3779}, {12'sd1250, 11'sd-906, 13'sd-3902}},
{{10'sd497, 13'sd-2703, 13'sd-4025}, {12'sd-1476, 10'sd381, 10'sd-286}, {13'sd-2321, 12'sd1343, 12'sd1210}},
{{13'sd-2248, 13'sd-3221, 1'sd0}, {13'sd-3877, 11'sd586, 11'sd-733}, {10'sd-446, 13'sd-2450, 13'sd3431}},
{{12'sd1700, 12'sd2038, 10'sd403}, {13'sd-2635, 12'sd1558, 13'sd2101}, {12'sd1644, 11'sd-747, 12'sd-1688}},
{{9'sd155, 10'sd508, 11'sd-845}, {12'sd1236, 13'sd2230, 8'sd106}, {12'sd-1332, 13'sd2382, 8'sd66}},
{{13'sd3420, 13'sd2941, 12'sd-1260}, {13'sd3879, 10'sd-493, 12'sd1595}, {13'sd2549, 12'sd1675, 13'sd-2817}},
{{11'sd-557, 12'sd-1247, 13'sd-2404}, {12'sd1369, 11'sd575, 8'sd-117}, {13'sd2675, 13'sd2384, 12'sd-1757}},
{{12'sd1436, 9'sd224, 13'sd3060}, {12'sd-1311, 12'sd1692, 12'sd1668}, {10'sd-441, 10'sd499, 12'sd-1941}},
{{10'sd-478, 12'sd1945, 11'sd-890}, {11'sd870, 13'sd2152, 13'sd-2762}, {13'sd-2277, 9'sd-233, 12'sd-1681}},
{{11'sd1000, 13'sd-2396, 11'sd-547}, {1'sd0, 13'sd-2823, 9'sd-206}, {11'sd-587, 11'sd-849, 13'sd2439}},
{{13'sd-3072, 12'sd-1541, 12'sd1137}, {13'sd-2128, 13'sd-2513, 11'sd-573}, {12'sd-1710, 11'sd-756, 8'sd115}},
{{12'sd-1031, 7'sd44, 12'sd-1904}, {12'sd1399, 11'sd-996, 10'sd-348}, {13'sd3096, 11'sd-753, 13'sd2160}},
{{10'sd467, 9'sd234, 11'sd828}, {12'sd1511, 9'sd227, 11'sd859}, {11'sd866, 9'sd-169, 12'sd1510}},
{{13'sd-2091, 12'sd1159, 12'sd1164}, {12'sd1087, 12'sd-1633, 12'sd1987}, {13'sd-3014, 11'sd873, 13'sd-2476}},
{{13'sd2951, 12'sd-1979, 9'sd213}, {13'sd3039, 11'sd-813, 13'sd-2629}, {11'sd612, 11'sd-991, 11'sd736}},
{{11'sd985, 10'sd-506, 13'sd2659}, {10'sd-436, 11'sd669, 12'sd-1714}, {11'sd634, 8'sd71, 12'sd1029}},
{{10'sd-367, 11'sd600, 13'sd-2057}, {12'sd-1259, 8'sd109, 12'sd1398}, {12'sd-1653, 13'sd-2454, 13'sd-2649}},
{{12'sd-1698, 12'sd-1837, 12'sd-1623}, {13'sd-2573, 12'sd-1965, 11'sd-560}, {13'sd-2260, 11'sd570, 12'sd-1411}},
{{13'sd-3969, 12'sd1089, 12'sd1761}, {12'sd-1874, 13'sd2093, 13'sd4070}, {13'sd-2094, 8'sd123, 13'sd3947}},
{{11'sd802, 11'sd750, 13'sd-2838}, {12'sd-1136, 13'sd2894, 13'sd-3460}, {13'sd-2393, 13'sd3162, 12'sd-1877}},
{{12'sd-1608, 11'sd802, 10'sd-352}, {9'sd135, 10'sd470, 12'sd1425}, {11'sd628, 11'sd-581, 13'sd2866}},
{{13'sd2563, 12'sd-1507, 10'sd421}, {8'sd88, 11'sd825, 12'sd1598}, {12'sd1711, 12'sd-1272, 12'sd-1771}},
{{11'sd-1006, 2'sd-1, 13'sd3591}, {12'sd1290, 9'sd215, 13'sd2731}, {13'sd-2118, 12'sd1702, 13'sd-2131}},
{{7'sd50, 11'sd944, 8'sd88}, {11'sd852, 13'sd2168, 13'sd-2123}, {12'sd-1968, 13'sd2406, 12'sd1747}},
{{13'sd3261, 8'sd-97, 13'sd2539}, {13'sd2601, 11'sd923, 10'sd379}, {13'sd4032, 11'sd959, 13'sd-2278}},
{{13'sd-2304, 6'sd-27, 12'sd-1864}, {13'sd-2228, 11'sd-730, 11'sd697}, {13'sd-2239, 13'sd2403, 12'sd-2031}},
{{13'sd-2780, 6'sd28, 7'sd47}, {12'sd-1366, 10'sd-434, 12'sd-1756}, {13'sd-2235, 13'sd-2995, 12'sd1822}},
{{12'sd-1602, 11'sd702, 12'sd-1972}, {11'sd807, 10'sd-285, 12'sd1718}, {13'sd-3837, 10'sd-443, 13'sd3095}},
{{13'sd2167, 13'sd-2518, 13'sd-2055}, {11'sd646, 12'sd1823, 12'sd1905}, {11'sd-708, 12'sd1150, 13'sd-3027}},
{{11'sd-710, 13'sd2227, 13'sd2235}, {12'sd1778, 13'sd-2658, 13'sd2996}, {11'sd-561, 12'sd-1319, 13'sd2117}},
{{7'sd-50, 12'sd-1976, 12'sd-1764}, {12'sd1451, 13'sd2147, 10'sd422}, {11'sd988, 13'sd-2244, 8'sd-120}},
{{12'sd-1578, 12'sd-1801, 11'sd-792}, {9'sd-160, 12'sd1268, 13'sd2495}, {11'sd-779, 13'sd2123, 12'sd1779}},
{{7'sd48, 12'sd-1616, 12'sd-1679}, {12'sd-1204, 11'sd864, 13'sd2343}, {11'sd-731, 13'sd2092, 7'sd63}},
{{12'sd-1253, 6'sd26, 13'sd2980}, {10'sd-477, 13'sd-2155, 12'sd-1082}, {9'sd215, 13'sd-2198, 11'sd744}},
{{9'sd174, 11'sd1010, 12'sd-1662}, {13'sd2425, 13'sd-2186, 12'sd-1595}, {13'sd-2406, 13'sd2944, 12'sd-1703}},
{{13'sd-2698, 13'sd2319, 12'sd-1901}, {13'sd2107, 9'sd225, 12'sd-1064}, {10'sd392, 11'sd744, 13'sd2091}},
{{13'sd2479, 11'sd765, 10'sd-468}, {11'sd882, 9'sd226, 9'sd-251}, {13'sd2583, 12'sd1380, 13'sd-2677}},
{{9'sd143, 12'sd1536, 12'sd1117}, {10'sd268, 10'sd494, 12'sd-1255}, {12'sd-1162, 12'sd1221, 11'sd-1004}},
{{14'sd5107, 11'sd-687, 13'sd-2535}, {11'sd905, 12'sd1044, 13'sd-2190}, {13'sd2448, 13'sd2580, 12'sd1450}},
{{8'sd120, 13'sd2649, 9'sd150}, {10'sd-494, 14'sd4256, 12'sd-1570}, {10'sd457, 13'sd2220, 10'sd-266}},
{{10'sd281, 12'sd1530, 13'sd2502}, {11'sd-899, 11'sd-710, 12'sd1637}, {10'sd347, 11'sd527, 12'sd-1815}},
{{12'sd-1188, 11'sd-764, 13'sd-2188}, {12'sd1804, 9'sd160, 10'sd-256}, {13'sd-2629, 12'sd-1442, 13'sd-2970}},
{{12'sd1852, 13'sd-2198, 12'sd1038}, {12'sd-1883, 9'sd201, 13'sd2193}, {12'sd-1855, 12'sd1527, 13'sd2519}},
{{12'sd1832, 8'sd83, 12'sd-1350}, {13'sd2333, 12'sd-1339, 13'sd-3689}, {12'sd-1690, 12'sd1465, 11'sd-710}},
{{13'sd3079, 11'sd-807, 13'sd3794}, {11'sd-629, 11'sd612, 12'sd1442}, {11'sd850, 7'sd-52, 11'sd-734}}},
{
{{13'sd-2502, 13'sd-3497, 12'sd-1974}, {11'sd981, 13'sd-3257, 9'sd162}, {12'sd1832, 12'sd-1100, 12'sd1377}},
{{11'sd1012, 12'sd-1615, 11'sd958}, {9'sd-183, 12'sd-1820, 12'sd1493}, {10'sd410, 12'sd-1821, 11'sd668}},
{{11'sd1023, 11'sd-853, 10'sd-459}, {13'sd-2661, 13'sd-2948, 10'sd-439}, {11'sd-778, 13'sd-2585, 11'sd-1015}},
{{12'sd1757, 13'sd-2627, 12'sd-1670}, {11'sd743, 8'sd102, 13'sd-2906}, {12'sd-1910, 12'sd-1569, 13'sd2456}},
{{9'sd193, 13'sd-2403, 9'sd205}, {9'sd-150, 9'sd-202, 12'sd1112}, {10'sd477, 13'sd-2237, 8'sd-94}},
{{11'sd970, 9'sd226, 12'sd-1667}, {10'sd-391, 12'sd1247, 13'sd2319}, {13'sd2781, 12'sd1208, 13'sd-2329}},
{{12'sd-1412, 11'sd-886, 13'sd2589}, {12'sd1697, 12'sd-1987, 13'sd-2121}, {12'sd-1667, 12'sd-1294, 13'sd-2259}},
{{11'sd-992, 13'sd2576, 12'sd1903}, {12'sd-1501, 11'sd756, 13'sd-2913}, {12'sd-1451, 12'sd-1048, 12'sd-1518}},
{{12'sd1422, 13'sd2170, 10'sd-274}, {12'sd-1643, 13'sd-2205, 12'sd1440}, {11'sd-815, 13'sd-2196, 13'sd2280}},
{{12'sd1395, 13'sd-2869, 13'sd-2305}, {10'sd-502, 12'sd1823, 12'sd-1508}, {11'sd-568, 11'sd690, 8'sd-111}},
{{9'sd-130, 11'sd705, 13'sd-3390}, {12'sd1407, 12'sd-1537, 13'sd-3735}, {12'sd-1133, 12'sd1071, 11'sd-756}},
{{13'sd-2544, 9'sd-223, 9'sd-129}, {9'sd144, 11'sd-608, 13'sd2635}, {13'sd2745, 12'sd1379, 13'sd-2129}},
{{12'sd-1853, 12'sd1147, 12'sd1541}, {10'sd-293, 11'sd-865, 11'sd-968}, {11'sd-540, 12'sd1757, 8'sd102}},
{{11'sd659, 13'sd-2182, 13'sd2732}, {13'sd-2340, 12'sd-1265, 12'sd1453}, {12'sd1044, 11'sd-683, 8'sd100}},
{{12'sd-1764, 13'sd-2323, 12'sd-1129}, {10'sd422, 12'sd1083, 12'sd1938}, {10'sd419, 12'sd1734, 12'sd2039}},
{{12'sd2022, 11'sd604, 13'sd2741}, {13'sd2324, 12'sd1480, 11'sd-737}, {13'sd2976, 11'sd-844, 11'sd-892}},
{{9'sd-190, 11'sd1018, 13'sd3099}, {13'sd-3057, 13'sd-3135, 11'sd842}, {8'sd-119, 13'sd-2211, 11'sd-617}},
{{12'sd1362, 13'sd-3601, 9'sd224}, {12'sd-1891, 13'sd-2234, 13'sd2291}, {13'sd2588, 14'sd-4140, 9'sd167}},
{{11'sd-859, 13'sd2506, 9'sd-216}, {12'sd-1942, 13'sd-2445, 10'sd-361}, {13'sd-2059, 8'sd-123, 13'sd2631}},
{{11'sd732, 13'sd-2235, 12'sd1071}, {11'sd-543, 12'sd-1320, 12'sd-2026}, {11'sd967, 11'sd-530, 12'sd-1478}},
{{11'sd768, 12'sd-1703, 11'sd-581}, {11'sd-831, 12'sd-1434, 13'sd2227}, {7'sd41, 13'sd2523, 13'sd-2542}},
{{13'sd2868, 12'sd1798, 13'sd-2165}, {12'sd1110, 12'sd1617, 12'sd-1210}, {9'sd-255, 12'sd1700, 8'sd-125}},
{{11'sd667, 12'sd-1107, 10'sd-363}, {13'sd-2235, 13'sd2345, 12'sd-1526}, {9'sd149, 12'sd-1639, 12'sd1296}},
{{12'sd-1318, 12'sd1611, 10'sd454}, {11'sd595, 11'sd526, 11'sd-728}, {12'sd1463, 12'sd1940, 10'sd475}},
{{11'sd1021, 13'sd-2782, 13'sd-2264}, {12'sd1946, 11'sd-919, 12'sd1327}, {13'sd3230, 11'sd583, 13'sd3050}},
{{12'sd1550, 13'sd2210, 12'sd-1445}, {10'sd-481, 13'sd2596, 11'sd-814}, {13'sd2930, 12'sd1248, 12'sd1927}},
{{12'sd-1943, 9'sd202, 12'sd-1333}, {12'sd-1358, 12'sd1996, 13'sd-2360}, {12'sd1333, 11'sd916, 12'sd-1899}},
{{11'sd545, 12'sd-1595, 13'sd2834}, {12'sd-1807, 11'sd953, 13'sd2086}, {13'sd2460, 12'sd1882, 12'sd-1219}},
{{12'sd1502, 6'sd-16, 11'sd-568}, {13'sd-2410, 13'sd2237, 11'sd-563}, {13'sd-3098, 13'sd-2178, 13'sd-2549}},
{{12'sd1169, 13'sd-2581, 12'sd1167}, {13'sd-2397, 13'sd2098, 11'sd-605}, {13'sd-3432, 11'sd-600, 13'sd-2278}},
{{12'sd2046, 10'sd-438, 9'sd198}, {13'sd2456, 12'sd1467, 13'sd-2605}, {11'sd831, 11'sd892, 11'sd-601}},
{{9'sd158, 13'sd-2490, 9'sd-227}, {13'sd-2247, 10'sd-289, 10'sd423}, {10'sd457, 13'sd-2402, 13'sd-2757}},
{{10'sd-496, 12'sd1874, 13'sd-2158}, {13'sd2234, 11'sd681, 11'sd1015}, {11'sd944, 11'sd-744, 11'sd-865}},
{{13'sd-2816, 13'sd2176, 12'sd-1949}, {11'sd793, 13'sd3052, 12'sd-1396}, {13'sd-2398, 12'sd1250, 13'sd-2163}},
{{12'sd1240, 13'sd2503, 11'sd813}, {13'sd-2444, 9'sd159, 11'sd-659}, {9'sd-206, 13'sd2925, 10'sd409}},
{{12'sd1836, 11'sd-881, 12'sd-1133}, {12'sd1842, 8'sd-124, 11'sd-578}, {13'sd-2118, 13'sd-2200, 13'sd2478}},
{{12'sd-2013, 12'sd1049, 12'sd1993}, {12'sd-1862, 10'sd-439, 11'sd952}, {13'sd-2836, 8'sd-122, 11'sd-937}},
{{12'sd1424, 13'sd-2362, 2'sd-1}, {12'sd1352, 10'sd370, 11'sd-869}, {12'sd-1060, 7'sd-45, 10'sd-351}},
{{12'sd1714, 12'sd1037, 11'sd522}, {11'sd-589, 6'sd-19, 6'sd-28}, {12'sd-1992, 12'sd-2047, 13'sd-2197}},
{{11'sd-637, 10'sd441, 9'sd247}, {12'sd1300, 12'sd1828, 12'sd1153}, {12'sd1879, 12'sd-1500, 13'sd-2439}},
{{13'sd-2190, 7'sd41, 11'sd711}, {13'sd2079, 9'sd219, 12'sd1369}, {12'sd1409, 11'sd766, 12'sd1391}},
{{10'sd261, 12'sd1511, 12'sd1440}, {8'sd-81, 13'sd-2083, 10'sd482}, {7'sd61, 12'sd-1194, 8'sd-65}},
{{11'sd655, 13'sd-2219, 13'sd-2500}, {12'sd-2016, 11'sd-759, 11'sd-606}, {12'sd1664, 12'sd1945, 12'sd-1368}},
{{11'sd-885, 13'sd2218, 8'sd-74}, {13'sd2357, 11'sd959, 12'sd-1143}, {11'sd650, 13'sd3436, 12'sd1232}},
{{13'sd2082, 10'sd-493, 13'sd2415}, {9'sd-217, 12'sd1314, 12'sd1889}, {12'sd1479, 13'sd2178, 7'sd45}},
{{10'sd354, 13'sd2262, 12'sd-1177}, {12'sd1954, 10'sd395, 12'sd1844}, {12'sd-1594, 13'sd-2156, 13'sd2134}},
{{12'sd1103, 10'sd437, 12'sd-1615}, {12'sd-1336, 13'sd2108, 13'sd2473}, {12'sd1587, 13'sd-3207, 12'sd1089}},
{{12'sd1709, 11'sd872, 13'sd-2477}, {11'sd-765, 10'sd-326, 8'sd81}, {12'sd1491, 13'sd2399, 11'sd-913}},
{{12'sd1509, 13'sd2582, 13'sd-2346}, {13'sd-2438, 11'sd-992, 12'sd-1482}, {12'sd-1889, 12'sd-1420, 10'sd338}},
{{10'sd506, 8'sd-73, 10'sd-348}, {12'sd1346, 12'sd-1757, 12'sd-1607}, {11'sd-747, 12'sd1235, 13'sd2072}},
{{12'sd1033, 13'sd2367, 11'sd-710}, {13'sd-2259, 13'sd-2149, 12'sd1509}, {12'sd-1487, 8'sd-72, 13'sd-2507}},
{{13'sd-2553, 11'sd-556, 13'sd2402}, {6'sd-22, 11'sd871, 12'sd1346}, {13'sd-2057, 11'sd871, 12'sd1966}},
{{13'sd3475, 13'sd3109, 13'sd2200}, {12'sd1360, 12'sd1620, 13'sd-2369}, {13'sd-3513, 13'sd-3297, 10'sd-328}},
{{7'sd-54, 11'sd-781, 12'sd-1262}, {11'sd-590, 11'sd783, 12'sd-1658}, {12'sd-1753, 12'sd1058, 9'sd-159}},
{{12'sd1839, 12'sd1724, 11'sd855}, {12'sd1293, 13'sd-2623, 12'sd-1842}, {6'sd25, 13'sd2113, 11'sd589}},
{{11'sd-738, 12'sd-1415, 13'sd-2255}, {12'sd-1341, 12'sd-1661, 12'sd1160}, {11'sd-567, 12'sd1749, 9'sd-240}},
{{11'sd969, 13'sd2524, 12'sd1143}, {9'sd-233, 10'sd-501, 12'sd1823}, {13'sd-2253, 11'sd-930, 11'sd-644}},
{{13'sd3142, 13'sd-3283, 12'sd2007}, {12'sd-1080, 13'sd-2747, 13'sd-2530}, {11'sd570, 13'sd2856, 10'sd414}},
{{11'sd668, 13'sd-2159, 12'sd1239}, {13'sd2620, 11'sd-758, 12'sd1572}, {12'sd1463, 13'sd2591, 11'sd-874}},
{{13'sd2321, 12'sd1560, 12'sd-1432}, {11'sd760, 9'sd237, 11'sd-1020}, {12'sd1902, 13'sd2453, 11'sd-565}},
{{12'sd1720, 11'sd951, 11'sd-929}, {8'sd90, 12'sd-1810, 12'sd1580}, {12'sd1764, 12'sd1589, 13'sd2207}},
{{11'sd-555, 11'sd-988, 12'sd-1896}, {13'sd2521, 10'sd-454, 11'sd-754}, {10'sd487, 11'sd818, 10'sd-485}},
{{11'sd-773, 12'sd1499, 11'sd-628}, {13'sd-2843, 13'sd-2531, 12'sd-1322}, {10'sd307, 9'sd178, 6'sd-27}},
{{12'sd-2037, 12'sd-1600, 12'sd1352}, {11'sd936, 13'sd2424, 12'sd-1659}, {11'sd526, 13'sd2542, 9'sd-134}}},
{
{{10'sd-328, 11'sd1009, 10'sd-348}, {12'sd-1526, 12'sd-1072, 6'sd-25}, {12'sd1281, 12'sd-1894, 10'sd379}},
{{10'sd435, 13'sd2579, 10'sd273}, {11'sd-978, 13'sd-2379, 12'sd-1166}, {12'sd-1580, 13'sd-2113, 11'sd629}},
{{12'sd1235, 12'sd-1356, 12'sd-1057}, {13'sd2102, 11'sd1017, 12'sd1186}, {13'sd2733, 13'sd2462, 10'sd-380}},
{{13'sd-2270, 13'sd2484, 10'sd443}, {11'sd867, 10'sd469, 11'sd543}, {12'sd1026, 12'sd1415, 12'sd1083}},
{{13'sd2064, 13'sd-2433, 13'sd-2866}, {9'sd178, 12'sd1858, 7'sd32}, {11'sd-580, 12'sd-1456, 13'sd-2930}},
{{12'sd1235, 13'sd-2101, 13'sd2754}, {10'sd485, 12'sd-1199, 13'sd-2502}, {12'sd-1248, 8'sd-95, 13'sd2135}},
{{12'sd1116, 10'sd342, 12'sd-1226}, {12'sd1630, 12'sd1314, 11'sd815}, {11'sd757, 13'sd-2576, 13'sd2220}},
{{11'sd766, 13'sd2280, 9'sd-166}, {12'sd1223, 13'sd-2829, 12'sd1430}, {12'sd1084, 12'sd-1694, 11'sd973}},
{{10'sd397, 12'sd1436, 12'sd1957}, {12'sd-1068, 13'sd-2396, 10'sd-378}, {12'sd-1881, 12'sd-1104, 11'sd-895}},
{{13'sd2272, 12'sd1789, 9'sd240}, {12'sd-1268, 12'sd-1692, 12'sd-1554}, {12'sd-1392, 12'sd-1814, 9'sd-130}},
{{14'sd4687, 13'sd3254, 11'sd911}, {14'sd5290, 13'sd2083, 13'sd2208}, {13'sd4051, 13'sd2797, 11'sd778}},
{{9'sd202, 12'sd-1769, 10'sd457}, {12'sd-1046, 12'sd1328, 11'sd562}, {10'sd-424, 11'sd-979, 12'sd-1786}},
{{12'sd1277, 13'sd2055, 12'sd1993}, {12'sd-1892, 13'sd-2301, 12'sd1204}, {11'sd717, 12'sd-1401, 9'sd138}},
{{12'sd1827, 12'sd1215, 13'sd2293}, {8'sd-126, 11'sd937, 13'sd-2271}, {11'sd938, 10'sd394, 11'sd690}},
{{11'sd727, 13'sd-2170, 12'sd-1319}, {12'sd1495, 10'sd-348, 13'sd2646}, {12'sd1378, 12'sd1680, 11'sd954}},
{{12'sd1810, 12'sd-1656, 12'sd-1103}, {12'sd1094, 13'sd2501, 11'sd-769}, {12'sd-1390, 9'sd176, 11'sd820}},
{{6'sd-25, 10'sd387, 12'sd1476}, {8'sd65, 12'sd-1286, 12'sd1047}, {13'sd-2730, 13'sd-2101, 12'sd1392}},
{{12'sd-1518, 11'sd514, 11'sd668}, {10'sd-421, 13'sd2679, 10'sd382}, {10'sd494, 13'sd3443, 12'sd2010}},
{{6'sd16, 12'sd1231, 11'sd650}, {12'sd1679, 10'sd-314, 12'sd1519}, {12'sd1982, 12'sd-1738, 8'sd-123}},
{{12'sd1413, 13'sd2702, 12'sd-1408}, {10'sd-465, 7'sd42, 11'sd-558}, {9'sd-157, 13'sd2477, 12'sd-1716}},
{{12'sd1116, 12'sd1839, 10'sd336}, {13'sd-2433, 12'sd-1771, 13'sd-2411}, {12'sd2025, 12'sd1613, 12'sd1581}},
{{12'sd1512, 12'sd1809, 11'sd777}, {12'sd-1892, 12'sd-1429, 9'sd187}, {12'sd1475, 13'sd-2305, 11'sd-555}},
{{12'sd-1341, 12'sd-1256, 13'sd-2324}, {13'sd2653, 13'sd2297, 11'sd911}, {12'sd-1980, 11'sd785, 11'sd-650}},
{{12'sd1699, 13'sd-2214, 13'sd-2800}, {12'sd-1877, 12'sd1479, 11'sd659}, {13'sd2514, 13'sd2792, 11'sd-597}},
{{14'sd-4472, 11'sd-834, 10'sd-372}, {13'sd-2075, 10'sd-326, 12'sd1690}, {11'sd-599, 12'sd-1348, 11'sd906}},
{{11'sd-916, 10'sd388, 13'sd2401}, {8'sd-124, 11'sd774, 12'sd1464}, {12'sd1731, 10'sd387, 12'sd1995}},
{{11'sd-755, 12'sd1472, 11'sd792}, {13'sd-2398, 12'sd1239, 12'sd-1657}, {12'sd1154, 12'sd1810, 12'sd-1378}},
{{12'sd1405, 11'sd-936, 12'sd-1511}, {9'sd244, 13'sd-2239, 12'sd1637}, {12'sd-1573, 13'sd2335, 12'sd-1217}},
{{12'sd-1507, 9'sd128, 11'sd-748}, {12'sd-2027, 12'sd2006, 12'sd1893}, {12'sd-1371, 5'sd9, 13'sd-2303}},
{{11'sd770, 12'sd1394, 13'sd-3069}, {10'sd372, 13'sd-2423, 11'sd-884}, {12'sd1833, 12'sd1587, 12'sd-1796}},
{{12'sd-1178, 13'sd2387, 12'sd1207}, {13'sd2524, 12'sd-1924, 12'sd-1097}, {10'sd495, 10'sd488, 8'sd-66}},
{{11'sd-572, 11'sd645, 8'sd126}, {9'sd-183, 12'sd1639, 12'sd1234}, {13'sd2648, 12'sd-1617, 4'sd7}},
{{12'sd1098, 13'sd2363, 12'sd-1980}, {8'sd-75, 13'sd-2132, 12'sd-1041}, {11'sd838, 12'sd1651, 13'sd2845}},
{{11'sd-812, 11'sd-623, 13'sd2291}, {12'sd1367, 12'sd-1967, 9'sd-226}, {12'sd-1224, 12'sd-1194, 13'sd2455}},
{{13'sd2615, 11'sd-814, 11'sd-1012}, {11'sd-916, 11'sd-673, 12'sd-1903}, {11'sd-519, 11'sd714, 12'sd1900}},
{{12'sd-1170, 10'sd-267, 10'sd-499}, {13'sd2434, 11'sd975, 12'sd1262}, {10'sd-471, 13'sd-2581, 10'sd-329}},
{{12'sd1319, 11'sd-718, 12'sd1753}, {11'sd-1002, 13'sd-2141, 12'sd-1705}, {12'sd1357, 11'sd-933, 11'sd906}},
{{9'sd-151, 8'sd-73, 12'sd-1968}, {13'sd-3550, 10'sd-360, 13'sd-2668}, {12'sd-2035, 13'sd-3023, 13'sd-3372}},
{{10'sd295, 11'sd684, 9'sd216}, {11'sd594, 12'sd1874, 13'sd2059}, {6'sd-23, 9'sd166, 13'sd-2209}},
{{12'sd1852, 12'sd-1205, 10'sd-357}, {13'sd2804, 13'sd2280, 12'sd-1736}, {12'sd1732, 8'sd-86, 13'sd-2326}},
{{13'sd-2706, 1'sd0, 8'sd-115}, {13'sd-2050, 13'sd-2760, 12'sd-1843}, {13'sd2428, 10'sd-349, 11'sd-642}},
{{12'sd1885, 13'sd-2708, 13'sd-2319}, {12'sd-1660, 12'sd-1540, 12'sd-1579}, {12'sd1165, 12'sd-1547, 10'sd-282}},
{{12'sd1165, 13'sd2503, 10'sd476}, {12'sd1592, 6'sd-25, 11'sd606}, {12'sd1622, 13'sd2133, 11'sd-813}},
{{12'sd-1904, 12'sd-1330, 13'sd2310}, {12'sd-1045, 13'sd2295, 13'sd2141}, {12'sd1343, 11'sd-712, 11'sd755}},
{{10'sd-490, 13'sd-2333, 12'sd1247}, {12'sd-1500, 12'sd1364, 13'sd-2727}, {9'sd241, 13'sd-2209, 12'sd1705}},
{{11'sd-593, 11'sd-610, 13'sd-2780}, {12'sd1977, 8'sd69, 13'sd-2083}, {9'sd-171, 9'sd-229, 12'sd-1240}},
{{9'sd235, 13'sd-2331, 13'sd2718}, {12'sd1997, 12'sd-1160, 12'sd-1458}, {12'sd1121, 12'sd1979, 12'sd1148}},
{{12'sd1476, 13'sd2121, 11'sd519}, {11'sd1010, 10'sd421, 13'sd-2130}, {12'sd-1681, 8'sd-93, 7'sd58}},
{{12'sd1560, 13'sd2273, 11'sd907}, {12'sd-1251, 13'sd-2445, 11'sd-560}, {13'sd-2370, 11'sd919, 12'sd-1797}},
{{12'sd-1350, 11'sd-519, 12'sd-1152}, {12'sd1853, 11'sd889, 12'sd-1624}, {11'sd-987, 12'sd1065, 12'sd-1980}},
{{12'sd-1736, 12'sd1208, 10'sd352}, {11'sd822, 8'sd115, 12'sd1795}, {12'sd1228, 13'sd-3120, 12'sd1937}},
{{9'sd154, 11'sd-865, 12'sd1860}, {10'sd320, 12'sd-1945, 13'sd-2248}, {13'sd-2563, 10'sd269, 13'sd2346}},
{{9'sd178, 10'sd312, 7'sd-51}, {11'sd-682, 12'sd-1834, 12'sd1200}, {13'sd2360, 13'sd2087, 12'sd-1139}},
{{11'sd-1016, 12'sd-1431, 10'sd503}, {11'sd-649, 12'sd1629, 11'sd670}, {11'sd-688, 11'sd-686, 13'sd2108}},
{{12'sd-1913, 13'sd-2420, 9'sd-202}, {12'sd-1359, 11'sd516, 11'sd-663}, {12'sd-1409, 12'sd1932, 11'sd-675}},
{{7'sd-63, 12'sd-1161, 11'sd-656}, {10'sd508, 12'sd-1681, 11'sd864}, {12'sd1520, 11'sd-946, 13'sd2469}},
{{8'sd-124, 10'sd-273, 11'sd924}, {9'sd-198, 11'sd-559, 9'sd-201}, {13'sd2672, 11'sd-524, 13'sd2904}},
{{11'sd810, 10'sd407, 11'sd540}, {11'sd-762, 13'sd-2693, 12'sd-1100}, {12'sd1658, 13'sd3247, 13'sd2529}},
{{10'sd483, 13'sd-3068, 13'sd-2473}, {11'sd-870, 12'sd1283, 9'sd-246}, {13'sd3576, 11'sd-753, 12'sd1033}},
{{11'sd-629, 12'sd-1779, 13'sd2078}, {13'sd2482, 12'sd-1590, 13'sd-2237}, {8'sd-114, 12'sd1794, 13'sd2239}},
{{13'sd-2210, 10'sd421, 12'sd1101}, {11'sd869, 11'sd929, 12'sd1887}, {12'sd-1104, 13'sd-2127, 13'sd-2109}},
{{10'sd-287, 12'sd-1571, 10'sd412}, {12'sd1403, 12'sd1559, 13'sd2049}, {12'sd-1577, 11'sd-699, 11'sd824}},
{{12'sd-1751, 13'sd-2586, 11'sd-631}, {11'sd921, 13'sd-2165, 13'sd2437}, {12'sd1224, 12'sd2045, 10'sd-359}},
{{13'sd-3757, 12'sd1970, 12'sd-1732}, {13'sd-3240, 12'sd-1615, 12'sd2031}, {12'sd-1288, 13'sd-2776, 11'sd763}}},
{
{{12'sd-1999, 12'sd-1077, 12'sd-1628}, {7'sd52, 13'sd-2859, 13'sd-3745}, {12'sd1168, 13'sd2302, 12'sd1086}},
{{11'sd-745, 12'sd-1033, 11'sd-864}, {13'sd2105, 12'sd1828, 11'sd785}, {12'sd1376, 10'sd-402, 13'sd-2320}},
{{13'sd3174, 11'sd-789, 12'sd-1641}, {7'sd49, 11'sd539, 12'sd-1792}, {12'sd-2042, 11'sd-866, 12'sd-1676}},
{{13'sd3144, 12'sd1754, 12'sd-1276}, {12'sd-1928, 12'sd1258, 12'sd-1852}, {10'sd-282, 12'sd1973, 12'sd1192}},
{{13'sd2345, 12'sd-1186, 11'sd674}, {11'sd-948, 12'sd1507, 7'sd34}, {13'sd2395, 7'sd40, 13'sd-2232}},
{{11'sd666, 12'sd1720, 13'sd-2895}, {12'sd2032, 11'sd781, 12'sd-1885}, {12'sd-1172, 12'sd1432, 13'sd-2143}},
{{11'sd969, 13'sd2335, 13'sd3064}, {10'sd332, 10'sd413, 12'sd-1545}, {10'sd358, 12'sd1805, 13'sd-2535}},
{{6'sd20, 10'sd394, 11'sd-529}, {12'sd-1339, 13'sd2290, 12'sd1355}, {13'sd2275, 12'sd1882, 13'sd-2145}},
{{10'sd285, 12'sd-1578, 13'sd-2055}, {13'sd-3125, 13'sd-2390, 12'sd1435}, {13'sd2111, 11'sd912, 11'sd-958}},
{{12'sd-1651, 12'sd1459, 13'sd-2139}, {11'sd-820, 13'sd2258, 13'sd-2572}, {12'sd2002, 12'sd1209, 11'sd-984}},
{{11'sd-796, 12'sd1777, 13'sd2941}, {12'sd1825, 9'sd-135, 9'sd-171}, {13'sd-3161, 14'sd4255, 13'sd3917}},
{{12'sd1650, 8'sd-75, 12'sd-1723}, {12'sd1466, 9'sd150, 12'sd1927}, {10'sd501, 13'sd-2673, 13'sd2746}},
{{12'sd-1870, 12'sd-1082, 12'sd1623}, {12'sd-1602, 7'sd-52, 12'sd-1151}, {12'sd-1302, 12'sd-1437, 12'sd-1331}},
{{11'sd-796, 12'sd1410, 12'sd-1341}, {12'sd-1765, 13'sd-2530, 12'sd1830}, {10'sd-289, 11'sd-827, 12'sd-1274}},
{{11'sd907, 13'sd2132, 12'sd1339}, {12'sd-1126, 12'sd-1696, 11'sd-964}, {13'sd-2614, 12'sd1377, 12'sd1938}},
{{13'sd2684, 12'sd1101, 13'sd2514}, {11'sd525, 12'sd-1971, 7'sd49}, {13'sd2803, 11'sd-718, 10'sd-508}},
{{12'sd-1419, 13'sd2542, 12'sd-1795}, {12'sd2032, 10'sd-445, 10'sd464}, {12'sd1526, 13'sd2617, 10'sd-473}},
{{11'sd541, 6'sd26, 13'sd-3976}, {10'sd494, 11'sd767, 10'sd-347}, {13'sd-2174, 12'sd-1859, 10'sd-404}},
{{11'sd-766, 12'sd1265, 11'sd-1011}, {12'sd-1916, 12'sd1341, 10'sd440}, {12'sd-1639, 12'sd1144, 7'sd-41}},
{{12'sd-1628, 12'sd-1546, 10'sd-507}, {13'sd-2153, 12'sd1186, 12'sd1211}, {12'sd-1837, 12'sd-1952, 10'sd361}},
{{12'sd1555, 10'sd-378, 12'sd-1993}, {13'sd-2476, 13'sd-2788, 13'sd2495}, {12'sd1426, 12'sd-1189, 10'sd344}},
{{13'sd-3818, 10'sd-407, 11'sd671}, {13'sd-3062, 13'sd2151, 8'sd117}, {5'sd-15, 9'sd219, 12'sd-1376}},
{{13'sd-3073, 12'sd-1458, 12'sd1193}, {11'sd-848, 11'sd862, 11'sd-699}, {12'sd1460, 12'sd1747, 13'sd-2212}},
{{12'sd1532, 12'sd1558, 12'sd-1767}, {13'sd-2689, 11'sd600, 13'sd2078}, {12'sd1389, 12'sd1290, 12'sd1277}},
{{11'sd-851, 11'sd590, 13'sd-3553}, {10'sd304, 12'sd1147, 11'sd998}, {11'sd-989, 11'sd721, 10'sd-297}},
{{11'sd-641, 13'sd-2455, 12'sd-1792}, {12'sd-2015, 12'sd1523, 13'sd-2677}, {13'sd-2492, 12'sd1043, 13'sd2135}},
{{12'sd-1830, 13'sd3193, 11'sd535}, {8'sd-96, 12'sd1455, 12'sd1178}, {12'sd-1186, 10'sd-318, 11'sd1018}},
{{11'sd-981, 11'sd-804, 13'sd2402}, {12'sd1978, 13'sd2182, 12'sd-2017}, {12'sd1046, 12'sd-1401, 12'sd-1830}},
{{10'sd-359, 13'sd2776, 12'sd-1463}, {13'sd2107, 12'sd-1192, 10'sd-403}, {9'sd135, 13'sd2116, 12'sd-1405}},
{{12'sd-1458, 13'sd2634, 12'sd-1057}, {12'sd1634, 12'sd-1179, 13'sd2585}, {13'sd-2196, 11'sd810, 12'sd-1422}},
{{11'sd-960, 9'sd149, 10'sd-320}, {11'sd-966, 11'sd830, 13'sd-2192}, {13'sd-2939, 11'sd-779, 6'sd30}},
{{13'sd2509, 12'sd-1994, 13'sd-3537}, {13'sd3246, 13'sd-2402, 13'sd-3454}, {13'sd2325, 13'sd-2065, 6'sd-27}},
{{12'sd1589, 13'sd-2325, 11'sd642}, {11'sd-624, 12'sd1822, 11'sd625}, {13'sd2091, 12'sd-1939, 10'sd-409}},
{{13'sd-2652, 13'sd-2741, 11'sd-622}, {12'sd-1699, 9'sd223, 12'sd-1451}, {11'sd776, 11'sd-512, 12'sd-1497}},
{{13'sd2303, 10'sd504, 11'sd-807}, {11'sd-834, 9'sd-142, 13'sd2815}, {9'sd172, 12'sd-1535, 12'sd1469}},
{{11'sd-628, 11'sd-703, 10'sd-428}, {9'sd-155, 11'sd-854, 11'sd807}, {12'sd-1724, 12'sd-1675, 12'sd-1309}},
{{13'sd-2498, 12'sd-1489, 10'sd-391}, {13'sd-2706, 11'sd-599, 13'sd2835}, {12'sd1089, 11'sd1018, 12'sd1619}},
{{11'sd813, 11'sd-769, 12'sd1470}, {13'sd2488, 12'sd1795, 12'sd-1591}, {11'sd623, 12'sd1127, 13'sd-2747}},
{{13'sd3260, 11'sd-626, 12'sd1495}, {13'sd2812, 11'sd-751, 12'sd-1607}, {13'sd2405, 12'sd-1647, 11'sd514}},
{{11'sd729, 11'sd-861, 11'sd949}, {13'sd3367, 12'sd1330, 12'sd1421}, {12'sd1856, 13'sd-2515, 13'sd2238}},
{{11'sd830, 13'sd2307, 10'sd-434}, {9'sd213, 12'sd-1644, 10'sd-320}, {11'sd946, 11'sd682, 12'sd-1789}},
{{13'sd3415, 13'sd-2157, 12'sd1025}, {12'sd-1599, 11'sd-750, 11'sd761}, {13'sd3176, 10'sd445, 12'sd-1135}},
{{11'sd-909, 12'sd-1675, 11'sd-757}, {9'sd189, 12'sd-1030, 13'sd-2049}, {12'sd-1503, 9'sd196, 11'sd879}},
{{11'sd-521, 12'sd1909, 12'sd1490}, {11'sd-732, 12'sd-1487, 13'sd2236}, {13'sd-2565, 12'sd1744, 11'sd585}},
{{13'sd-3415, 11'sd847, 13'sd2347}, {10'sd432, 11'sd-732, 12'sd1940}, {9'sd-147, 13'sd2272, 13'sd-2941}},
{{10'sd-346, 12'sd-1745, 12'sd2005}, {8'sd85, 12'sd1460, 12'sd1192}, {12'sd1798, 12'sd-1165, 12'sd1732}},
{{13'sd3360, 13'sd-2135, 9'sd197}, {12'sd-1728, 11'sd713, 13'sd-2517}, {13'sd-2499, 11'sd-942, 12'sd-1452}},
{{11'sd-968, 12'sd-1618, 12'sd-1965}, {12'sd-1691, 10'sd-481, 11'sd994}, {10'sd346, 12'sd2030, 13'sd2523}},
{{11'sd619, 13'sd2180, 12'sd-2038}, {12'sd1852, 12'sd-1127, 7'sd34}, {12'sd1600, 12'sd-1508, 12'sd-1281}},
{{4'sd5, 12'sd1332, 10'sd-299}, {13'sd2321, 13'sd2359, 6'sd30}, {13'sd-2882, 13'sd-2694, 11'sd-631}},
{{12'sd1974, 13'sd-2317, 12'sd-1953}, {13'sd2440, 11'sd-956, 12'sd-1329}, {12'sd1280, 12'sd-1321, 12'sd1035}},
{{11'sd-736, 12'sd1829, 10'sd456}, {10'sd329, 13'sd-2412, 13'sd2709}, {9'sd166, 5'sd-12, 12'sd1954}},
{{12'sd1965, 12'sd-1643, 12'sd-1202}, {13'sd2103, 12'sd-1975, 9'sd-215}, {12'sd1814, 13'sd-2975, 7'sd60}},
{{11'sd564, 11'sd582, 12'sd-1458}, {13'sd2144, 13'sd-3129, 13'sd-2561}, {11'sd797, 13'sd-2890, 11'sd931}},
{{11'sd796, 12'sd1835, 10'sd421}, {8'sd79, 13'sd2253, 9'sd179}, {12'sd1606, 10'sd296, 13'sd2260}},
{{11'sd-584, 10'sd-285, 12'sd1208}, {11'sd-770, 10'sd309, 10'sd498}, {12'sd-1213, 12'sd1595, 12'sd-1711}},
{{11'sd-1022, 13'sd2144, 11'sd866}, {11'sd-873, 13'sd3112, 12'sd1868}, {12'sd1532, 13'sd-2436, 11'sd920}},
{{12'sd1037, 11'sd826, 13'sd-2427}, {11'sd692, 11'sd594, 13'sd-2639}, {9'sd-217, 10'sd-380, 12'sd1700}},
{{13'sd-2313, 12'sd1436, 12'sd-1907}, {13'sd2959, 12'sd1078, 13'sd-2650}, {12'sd1914, 13'sd-2398, 12'sd-1652}},
{{10'sd-269, 9'sd230, 11'sd-878}, {13'sd2612, 12'sd-1936, 12'sd1327}, {13'sd-2056, 11'sd-768, 12'sd1340}},
{{8'sd-104, 13'sd2566, 12'sd-1670}, {9'sd-225, 11'sd-536, 13'sd-2735}, {13'sd-2369, 12'sd1645, 13'sd-2483}},
{{13'sd2844, 11'sd-598, 13'sd3005}, {13'sd2203, 9'sd-140, 12'sd1606}, {12'sd-1512, 11'sd-979, 10'sd364}},
{{10'sd329, 12'sd1768, 13'sd-3175}, {12'sd-1677, 11'sd533, 9'sd238}, {11'sd611, 10'sd-399, 10'sd-300}},
{{11'sd-664, 12'sd1893, 5'sd13}, {9'sd219, 13'sd-2373, 12'sd1311}, {10'sd-453, 11'sd-648, 13'sd2324}}},
{
{{12'sd-1151, 12'sd-1533, 9'sd-180}, {13'sd2916, 8'sd115, 13'sd-2270}, {12'sd1928, 13'sd2371, 11'sd579}},
{{12'sd-1413, 11'sd990, 13'sd-2220}, {13'sd2270, 12'sd1460, 12'sd1142}, {11'sd798, 13'sd-3398, 11'sd857}},
{{13'sd2295, 12'sd-1432, 12'sd1319}, {14'sd4401, 10'sd-383, 11'sd608}, {9'sd170, 13'sd-2782, 12'sd-1171}},
{{13'sd-2224, 10'sd382, 13'sd-2114}, {11'sd-852, 12'sd1326, 11'sd-586}, {10'sd331, 12'sd-1111, 12'sd1881}},
{{10'sd-390, 13'sd3207, 11'sd-557}, {10'sd305, 13'sd4000, 8'sd-102}, {13'sd2156, 12'sd1242, 13'sd3613}},
{{9'sd190, 12'sd1760, 10'sd352}, {13'sd2082, 13'sd2134, 11'sd795}, {12'sd1639, 11'sd-512, 12'sd-1511}},
{{13'sd2441, 12'sd1213, 12'sd-1796}, {13'sd-2663, 12'sd-1352, 10'sd261}, {13'sd-3296, 12'sd-1102, 11'sd-910}},
{{12'sd1798, 11'sd845, 12'sd-1966}, {13'sd2073, 13'sd-2755, 13'sd-2593}, {14'sd7388, 14'sd5187, 12'sd1857}},
{{12'sd-1299, 11'sd-528, 13'sd-2357}, {11'sd-706, 12'sd1749, 12'sd1682}, {13'sd2684, 13'sd2131, 12'sd1734}},
{{13'sd2325, 13'sd2611, 14'sd4304}, {12'sd-1765, 11'sd982, 13'sd2447}, {11'sd749, 13'sd2234, 11'sd1019}},
{{13'sd3257, 12'sd1359, 10'sd-466}, {13'sd-2301, 12'sd1052, 11'sd-521}, {11'sd904, 12'sd1309, 14'sd4996}},
{{13'sd-3425, 13'sd-2641, 13'sd-2570}, {13'sd2319, 10'sd496, 13'sd3444}, {10'sd-429, 13'sd2903, 11'sd-529}},
{{13'sd-2667, 11'sd-732, 13'sd-2469}, {14'sd-4473, 14'sd-5534, 10'sd-387}, {10'sd-264, 13'sd-2405, 12'sd1332}},
{{11'sd-1022, 12'sd1180, 12'sd-1081}, {9'sd252, 10'sd284, 12'sd1961}, {11'sd735, 12'sd-1365, 13'sd3293}},
{{13'sd3465, 10'sd380, 13'sd2663}, {12'sd-1374, 9'sd181, 13'sd-2762}, {12'sd-1710, 11'sd-830, 12'sd1505}},
{{13'sd2669, 10'sd352, 12'sd-1156}, {10'sd-272, 12'sd2015, 13'sd-2926}, {13'sd3704, 5'sd-11, 12'sd1135}},
{{13'sd-3400, 13'sd-3943, 8'sd-123}, {11'sd-808, 11'sd881, 13'sd-2384}, {9'sd-240, 13'sd-3404, 10'sd388}},
{{14'sd4280, 13'sd2556, 13'sd3315}, {13'sd2230, 9'sd212, 11'sd-670}, {12'sd2007, 11'sd557, 10'sd309}},
{{9'sd-242, 10'sd277, 10'sd411}, {12'sd2026, 13'sd-2205, 11'sd588}, {3'sd-3, 12'sd-1893, 12'sd-1043}},
{{9'sd-231, 12'sd2023, 9'sd-165}, {8'sd-125, 13'sd2321, 10'sd-399}, {13'sd2151, 11'sd-923, 12'sd1979}},
{{13'sd-2350, 13'sd2826, 6'sd18}, {13'sd2953, 11'sd-987, 11'sd545}, {12'sd-1268, 12'sd1323, 11'sd-698}},
{{13'sd3476, 13'sd2664, 13'sd3068}, {13'sd-3773, 13'sd-3846, 9'sd-253}, {15'sd-8342, 14'sd-4421, 12'sd-1550}},
{{10'sd332, 13'sd2391, 12'sd-1448}, {11'sd839, 12'sd-1333, 12'sd-1383}, {10'sd385, 11'sd-630, 12'sd-1594}},
{{13'sd3439, 10'sd-356, 11'sd-995}, {9'sd-133, 13'sd2831, 10'sd343}, {12'sd1751, 13'sd2217, 12'sd-1095}},
{{11'sd-665, 12'sd-1821, 10'sd-267}, {13'sd2801, 11'sd633, 14'sd4534}, {11'sd1001, 14'sd-4114, 7'sd35}},
{{11'sd863, 12'sd-1238, 9'sd200}, {9'sd224, 11'sd836, 10'sd-294}, {13'sd-2364, 11'sd-617, 11'sd789}},
{{12'sd-1127, 13'sd-2141, 10'sd424}, {12'sd-1793, 12'sd-1550, 11'sd993}, {13'sd-2511, 13'sd3021, 12'sd-1201}},
{{11'sd835, 12'sd1218, 13'sd3296}, {10'sd-356, 13'sd2183, 12'sd1952}, {11'sd910, 9'sd-131, 13'sd3586}},
{{8'sd-100, 9'sd201, 10'sd-370}, {14'sd-4647, 13'sd-3086, 11'sd-699}, {13'sd-3104, 12'sd-1125, 13'sd2492}},
{{12'sd-1131, 12'sd1331, 12'sd1139}, {13'sd-3796, 12'sd-1084, 12'sd1748}, {13'sd-2960, 12'sd1647, 12'sd-1712}},
{{13'sd-2227, 11'sd649, 11'sd-820}, {12'sd1949, 12'sd2021, 12'sd1670}, {11'sd830, 13'sd-2432, 12'sd-1167}},
{{6'sd-16, 10'sd460, 12'sd-1923}, {10'sd440, 13'sd-2285, 13'sd-3169}, {13'sd3777, 12'sd1944, 12'sd1092}},
{{11'sd656, 10'sd373, 11'sd957}, {12'sd1530, 11'sd-674, 12'sd-1076}, {10'sd-409, 13'sd-3824, 13'sd-2125}},
{{10'sd312, 13'sd-2238, 11'sd607}, {10'sd416, 11'sd588, 13'sd3410}, {10'sd-417, 12'sd1253, 12'sd1461}},
{{11'sd-737, 12'sd-1789, 13'sd-2941}, {11'sd514, 13'sd-2361, 13'sd-2478}, {11'sd682, 10'sd-416, 13'sd-2734}},
{{11'sd851, 12'sd-1911, 13'sd2193}, {12'sd1627, 12'sd1613, 13'sd2129}, {13'sd2078, 13'sd2697, 11'sd-625}},
{{12'sd1404, 12'sd-1307, 13'sd-2199}, {11'sd892, 10'sd-374, 13'sd2202}, {11'sd549, 13'sd2241, 11'sd671}},
{{11'sd725, 13'sd2169, 11'sd-539}, {8'sd-91, 13'sd-2507, 14'sd-4517}, {13'sd3500, 13'sd2316, 9'sd-142}},
{{12'sd-1778, 13'sd2058, 12'sd-1710}, {12'sd-1661, 12'sd1339, 11'sd567}, {13'sd-2709, 11'sd-1003, 12'sd1256}},
{{12'sd-1806, 13'sd-3232, 8'sd92}, {11'sd-1016, 12'sd-1433, 9'sd217}, {13'sd3068, 10'sd-443, 12'sd-1567}},
{{11'sd744, 12'sd-1912, 12'sd1143}, {11'sd-832, 9'sd-146, 12'sd-1983}, {11'sd-709, 13'sd-2150, 11'sd874}},
{{12'sd-1564, 12'sd1762, 10'sd463}, {13'sd-2301, 12'sd1978, 11'sd703}, {13'sd3193, 13'sd2117, 11'sd581}},
{{13'sd-2541, 9'sd-168, 13'sd-2395}, {12'sd-1438, 11'sd-674, 13'sd2502}, {13'sd3013, 9'sd255, 13'sd-2128}},
{{14'sd-4585, 10'sd344, 13'sd-3638}, {11'sd-721, 9'sd-248, 12'sd1961}, {10'sd-314, 13'sd3102, 13'sd2827}},
{{6'sd26, 12'sd1922, 12'sd-1663}, {13'sd-2399, 13'sd2543, 13'sd2438}, {12'sd1631, 12'sd-1650, 13'sd-2678}},
{{9'sd186, 13'sd3246, 13'sd2559}, {6'sd-31, 10'sd-333, 9'sd-147}, {12'sd1950, 12'sd-1717, 12'sd-1329}},
{{12'sd-2015, 13'sd-3087, 12'sd2002}, {13'sd-2917, 12'sd-1553, 10'sd267}, {13'sd-2771, 11'sd777, 11'sd667}},
{{5'sd10, 11'sd721, 11'sd-854}, {8'sd78, 12'sd-1615, 6'sd20}, {8'sd-125, 12'sd-1690, 11'sd-995}},
{{12'sd1067, 13'sd2234, 12'sd1357}, {12'sd-1776, 13'sd-2270, 12'sd-1464}, {8'sd92, 9'sd230, 13'sd2488}},
{{13'sd-2489, 11'sd-662, 12'sd1242}, {11'sd878, 10'sd-444, 12'sd-1745}, {12'sd1535, 13'sd-2773, 13'sd-2661}},
{{11'sd588, 9'sd243, 13'sd2647}, {13'sd-3090, 13'sd-2229, 10'sd-283}, {12'sd1276, 12'sd1444, 11'sd-602}},
{{8'sd-92, 12'sd1919, 10'sd-410}, {12'sd-1913, 12'sd1889, 12'sd1762}, {11'sd663, 12'sd-1142, 13'sd-2193}},
{{13'sd2965, 13'sd3252, 11'sd646}, {13'sd-2582, 13'sd-2313, 9'sd253}, {13'sd-3605, 13'sd-2917, 11'sd-816}},
{{13'sd3267, 11'sd769, 10'sd-417}, {10'sd421, 12'sd-1530, 13'sd-3004}, {11'sd772, 10'sd497, 12'sd-1085}},
{{13'sd2641, 12'sd-1720, 9'sd-248}, {13'sd3031, 12'sd-1850, 11'sd922}, {12'sd-1052, 13'sd-3444, 11'sd-540}},
{{12'sd1908, 12'sd-1364, 11'sd-922}, {13'sd2325, 13'sd-2488, 9'sd-224}, {12'sd2014, 12'sd1083, 10'sd-371}},
{{12'sd-1364, 13'sd2695, 12'sd-1085}, {12'sd-1029, 12'sd1756, 13'sd2856}, {11'sd-773, 12'sd1138, 13'sd-2994}},
{{13'sd2082, 12'sd1314, 13'sd-3899}, {12'sd-1440, 11'sd935, 13'sd-3836}, {7'sd53, 11'sd854, 11'sd-649}},
{{11'sd-538, 13'sd3648, 12'sd1583}, {11'sd521, 9'sd-167, 10'sd280}, {12'sd1300, 12'sd-1035, 11'sd1001}},
{{13'sd-2532, 12'sd-1201, 13'sd-2330}, {11'sd626, 13'sd-2359, 13'sd2700}, {11'sd827, 9'sd131, 11'sd-533}},
{{9'sd-236, 11'sd514, 8'sd-104}, {13'sd3076, 12'sd1991, 12'sd1382}, {11'sd867, 12'sd-1904, 13'sd-2060}},
{{12'sd-1094, 12'sd1870, 11'sd774}, {13'sd-2721, 12'sd1771, 11'sd761}, {12'sd1557, 10'sd416, 12'sd1300}},
{{12'sd-1423, 12'sd-1739, 11'sd543}, {12'sd1079, 8'sd-65, 12'sd1768}, {11'sd-707, 13'sd3079, 11'sd-546}},
{{12'sd1578, 12'sd1933, 12'sd1144}, {13'sd-2603, 13'sd2119, 12'sd1165}, {13'sd-2054, 12'sd-1151, 11'sd-740}}},
{
{{12'sd1152, 12'sd-2023, 13'sd2564}, {10'sd-435, 11'sd555, 13'sd2956}, {12'sd1242, 12'sd1218, 13'sd-2143}},
{{11'sd-854, 11'sd791, 11'sd-589}, {12'sd1556, 13'sd2540, 12'sd1307}, {10'sd443, 11'sd728, 13'sd2672}},
{{13'sd-2738, 9'sd186, 10'sd-491}, {13'sd2102, 10'sd-442, 11'sd-827}, {11'sd-757, 6'sd25, 10'sd299}},
{{11'sd-707, 11'sd766, 13'sd-2168}, {11'sd517, 12'sd1451, 13'sd-2451}, {12'sd1430, 10'sd477, 12'sd2037}},
{{12'sd1174, 8'sd-120, 12'sd-1959}, {12'sd-1967, 12'sd-1986, 13'sd2621}, {12'sd1566, 8'sd-73, 12'sd1944}},
{{13'sd2058, 12'sd1291, 12'sd1503}, {12'sd1048, 10'sd-493, 11'sd-620}, {13'sd2377, 12'sd-1505, 11'sd651}},
{{13'sd-2205, 12'sd-1212, 12'sd-1941}, {9'sd-239, 13'sd-2529, 13'sd-2436}, {11'sd-646, 12'sd-1413, 13'sd-2240}},
{{13'sd-2399, 11'sd-1023, 12'sd-1944}, {8'sd113, 11'sd-673, 13'sd2153}, {10'sd341, 13'sd-2075, 11'sd-626}},
{{12'sd1352, 11'sd543, 12'sd1259}, {10'sd485, 12'sd-1428, 13'sd2675}, {10'sd-465, 10'sd-465, 11'sd527}},
{{12'sd-2038, 11'sd735, 9'sd-191}, {12'sd-1735, 10'sd363, 12'sd-1613}, {9'sd-199, 11'sd843, 12'sd-1414}},
{{13'sd3867, 10'sd-438, 12'sd1986}, {8'sd72, 12'sd1195, 11'sd-715}, {11'sd-680, 10'sd420, 13'sd-3705}},
{{13'sd-2663, 13'sd2102, 12'sd-1422}, {12'sd-1807, 13'sd-2266, 12'sd1670}, {11'sd897, 10'sd-324, 12'sd1521}},
{{12'sd-1908, 12'sd-1814, 10'sd347}, {10'sd-481, 12'sd-1356, 13'sd2773}, {11'sd-939, 12'sd-1975, 13'sd-2182}},
{{13'sd2163, 13'sd2580, 12'sd1701}, {12'sd1396, 12'sd1985, 13'sd-2674}, {11'sd689, 13'sd2573, 11'sd-752}},
{{11'sd879, 12'sd-1252, 11'sd-934}, {11'sd-512, 11'sd-697, 13'sd-2510}, {12'sd1704, 9'sd-150, 10'sd-316}},
{{12'sd1787, 12'sd1403, 12'sd-1613}, {11'sd951, 13'sd2219, 11'sd-726}, {11'sd-684, 8'sd-66, 11'sd-612}},
{{10'sd423, 13'sd-2274, 12'sd1820}, {12'sd-1471, 13'sd-2443, 11'sd976}, {9'sd-237, 12'sd-1070, 12'sd-1823}},
{{14'sd-4458, 7'sd52, 10'sd-289}, {14'sd-4468, 13'sd-2466, 10'sd-285}, {12'sd1479, 12'sd-1345, 12'sd1700}},
{{10'sd-394, 13'sd-2767, 11'sd-662}, {12'sd1683, 11'sd-961, 12'sd1948}, {12'sd-2001, 12'sd-1696, 7'sd-33}},
{{11'sd1015, 11'sd881, 12'sd2006}, {12'sd1085, 11'sd-619, 12'sd1838}, {12'sd-2042, 12'sd-1143, 12'sd2017}},
{{11'sd563, 12'sd-1188, 11'sd-631}, {8'sd-67, 13'sd2661, 12'sd-1117}, {12'sd-1072, 13'sd-2655, 11'sd683}},
{{13'sd2300, 12'sd1363, 13'sd-2796}, {13'sd-2493, 12'sd2047, 12'sd1914}, {12'sd-1654, 12'sd1803, 10'sd-265}},
{{12'sd1463, 12'sd-1927, 11'sd533}, {8'sd116, 12'sd1734, 12'sd1658}, {12'sd1308, 12'sd-1391, 13'sd2381}},
{{9'sd-132, 12'sd-1512, 10'sd-337}, {13'sd2069, 13'sd2606, 12'sd-1873}, {10'sd-505, 11'sd875, 13'sd-2643}},
{{12'sd-1770, 11'sd616, 11'sd-516}, {13'sd-2732, 13'sd2128, 10'sd-464}, {12'sd1892, 13'sd2178, 12'sd-1565}},
{{12'sd-1748, 12'sd1226, 11'sd-554}, {9'sd132, 11'sd667, 13'sd2427}, {11'sd530, 10'sd-407, 12'sd1729}},
{{11'sd-998, 13'sd2413, 12'sd1798}, {13'sd2770, 11'sd581, 12'sd1333}, {9'sd-228, 12'sd-1380, 7'sd-43}},
{{12'sd-2039, 12'sd-1457, 12'sd-1987}, {11'sd-574, 13'sd2341, 12'sd1370}, {12'sd-1355, 9'sd-217, 11'sd-936}},
{{12'sd1410, 13'sd-2330, 12'sd1032}, {13'sd2559, 12'sd-1823, 11'sd-999}, {13'sd2453, 13'sd-2225, 12'sd1546}},
{{11'sd-643, 10'sd418, 10'sd-479}, {12'sd1565, 11'sd819, 12'sd1767}, {13'sd3015, 10'sd-398, 12'sd-1302}},
{{13'sd2751, 8'sd-68, 7'sd34}, {12'sd-2036, 11'sd-872, 11'sd632}, {12'sd-1574, 11'sd-702, 11'sd-702}},
{{10'sd432, 10'sd-335, 11'sd775}, {12'sd-2034, 10'sd289, 11'sd-698}, {11'sd804, 13'sd2057, 13'sd2269}},
{{13'sd2315, 11'sd977, 7'sd43}, {13'sd-2871, 12'sd-1604, 13'sd2205}, {10'sd386, 11'sd-746, 8'sd108}},
{{12'sd1900, 12'sd-1543, 13'sd2586}, {12'sd1272, 10'sd434, 11'sd-866}, {12'sd-1461, 10'sd-328, 10'sd450}},
{{9'sd228, 9'sd-210, 12'sd-2024}, {13'sd-2342, 13'sd-2377, 10'sd-274}, {11'sd995, 11'sd-543, 12'sd1492}},
{{13'sd2193, 12'sd1860, 11'sd-517}, {10'sd-418, 13'sd2789, 12'sd-1449}, {13'sd2271, 9'sd180, 13'sd-2720}},
{{8'sd-103, 13'sd2583, 11'sd796}, {9'sd201, 12'sd-1729, 13'sd-2555}, {12'sd1217, 11'sd789, 12'sd1221}},
{{10'sd377, 12'sd1813, 10'sd-420}, {11'sd-883, 10'sd-482, 12'sd1492}, {13'sd2622, 11'sd751, 13'sd2404}},
{{11'sd718, 13'sd-2254, 12'sd2022}, {9'sd-141, 10'sd454, 13'sd2544}, {12'sd1482, 11'sd810, 13'sd-2224}},
{{11'sd717, 10'sd-472, 12'sd1819}, {13'sd2523, 10'sd442, 11'sd-571}, {13'sd-2554, 13'sd2083, 12'sd-1319}},
{{9'sd194, 11'sd-1007, 13'sd3387}, {13'sd-2362, 11'sd851, 12'sd2004}, {12'sd-1913, 12'sd-1542, 12'sd1104}},
{{12'sd-1969, 11'sd610, 9'sd235}, {13'sd-2197, 12'sd-1635, 13'sd2596}, {12'sd1116, 12'sd1930, 12'sd-1838}},
{{12'sd-1188, 13'sd2571, 12'sd1545}, {9'sd-138, 13'sd-2101, 12'sd-1172}, {9'sd-249, 13'sd-2155, 11'sd839}},
{{9'sd-193, 13'sd2829, 12'sd-1773}, {12'sd1184, 9'sd-234, 12'sd-1468}, {12'sd-1204, 11'sd750, 13'sd-2316}},
{{13'sd2642, 12'sd1530, 13'sd-2146}, {10'sd-481, 12'sd-1504, 13'sd2412}, {11'sd624, 11'sd661, 12'sd1535}},
{{12'sd1428, 13'sd2312, 13'sd-2474}, {12'sd-2002, 12'sd-1071, 10'sd264}, {12'sd-1451, 13'sd-2054, 13'sd-2493}},
{{13'sd-2482, 11'sd752, 13'sd-2161}, {12'sd2033, 11'sd-633, 12'sd-1496}, {11'sd-1010, 13'sd3192, 11'sd1006}},
{{11'sd-513, 13'sd-2224, 11'sd623}, {12'sd1305, 11'sd946, 12'sd-1469}, {11'sd-743, 7'sd-62, 12'sd1969}},
{{13'sd-2476, 12'sd-1184, 11'sd-650}, {13'sd2629, 12'sd-1986, 13'sd-2749}, {12'sd1753, 12'sd1251, 10'sd304}},
{{12'sd-1993, 10'sd-347, 12'sd-1651}, {13'sd2563, 11'sd605, 13'sd2261}, {13'sd-2362, 10'sd456, 13'sd-2485}},
{{4'sd7, 11'sd692, 13'sd2477}, {13'sd2440, 11'sd560, 12'sd-2018}, {10'sd-496, 11'sd-717, 11'sd-731}},
{{12'sd-1531, 12'sd-1596, 10'sd415}, {11'sd-922, 12'sd1188, 12'sd-1192}, {12'sd-1238, 6'sd21, 12'sd1646}},
{{10'sd357, 12'sd1037, 11'sd660}, {13'sd-2173, 13'sd-2259, 12'sd-1996}, {13'sd2748, 11'sd583, 13'sd2450}},
{{12'sd-1209, 12'sd1549, 13'sd2591}, {12'sd-1604, 13'sd-2773, 11'sd905}, {12'sd-1475, 13'sd-2290, 12'sd-1281}},
{{13'sd-2098, 12'sd-1213, 13'sd2608}, {12'sd-1224, 13'sd-2753, 9'sd202}, {12'sd1374, 13'sd-2085, 13'sd-2456}},
{{11'sd-995, 11'sd515, 12'sd-1450}, {13'sd-2101, 10'sd-323, 11'sd-750}, {12'sd-1541, 13'sd2443, 13'sd2056}},
{{11'sd900, 5'sd-14, 11'sd699}, {12'sd-1325, 12'sd1238, 9'sd-213}, {12'sd1786, 12'sd1653, 10'sd323}},
{{7'sd46, 12'sd-1202, 10'sd279}, {9'sd172, 11'sd567, 12'sd-1222}, {11'sd812, 11'sd-876, 11'sd-935}},
{{12'sd-1961, 12'sd1731, 12'sd-1555}, {11'sd-922, 12'sd-1172, 12'sd1236}, {12'sd-1887, 12'sd1491, 13'sd3006}},
{{12'sd1613, 12'sd-1849, 12'sd1936}, {8'sd-126, 12'sd1910, 13'sd-2224}, {12'sd1333, 13'sd2367, 13'sd-2379}},
{{12'sd-1132, 11'sd585, 12'sd1803}, {13'sd2255, 13'sd2414, 12'sd-1962}, {12'sd1742, 9'sd-191, 12'sd1581}},
{{13'sd2530, 13'sd-2290, 12'sd1121}, {13'sd-2256, 10'sd-440, 11'sd843}, {11'sd834, 12'sd1977, 12'sd1203}},
{{13'sd-2704, 11'sd973, 13'sd3253}, {12'sd1334, 11'sd694, 12'sd1441}, {12'sd-1389, 11'sd-519, 13'sd2219}},
{{13'sd-3167, 11'sd984, 10'sd266}, {13'sd-2308, 13'sd2302, 13'sd2485}, {11'sd-623, 9'sd231, 12'sd1602}}},
{
{{8'sd-125, 10'sd-264, 12'sd1333}, {10'sd429, 12'sd-1175, 12'sd1370}, {12'sd-1778, 13'sd2491, 12'sd1710}},
{{12'sd1696, 13'sd-2554, 12'sd1191}, {11'sd-520, 13'sd-2688, 12'sd-1821}, {12'sd1613, 12'sd-1934, 12'sd1317}},
{{13'sd-3100, 13'sd-2346, 12'sd-1123}, {13'sd-2463, 7'sd-34, 12'sd1668}, {11'sd870, 12'sd1313, 11'sd888}},
{{9'sd248, 13'sd2545, 10'sd-480}, {11'sd876, 13'sd2461, 11'sd-728}, {10'sd-460, 12'sd1774, 11'sd-825}},
{{13'sd2181, 11'sd645, 12'sd-1895}, {13'sd-2592, 11'sd-635, 13'sd-2162}, {13'sd2178, 12'sd1626, 12'sd1470}},
{{12'sd-1592, 12'sd-1284, 10'sd-312}, {9'sd-196, 11'sd-828, 13'sd2701}, {13'sd2134, 12'sd-1717, 11'sd664}},
{{13'sd-2527, 13'sd-2590, 11'sd602}, {12'sd1223, 12'sd1154, 11'sd-677}, {12'sd-1653, 12'sd2021, 12'sd2005}},
{{13'sd2247, 13'sd3404, 13'sd-2419}, {9'sd-188, 11'sd-840, 12'sd1340}, {12'sd1753, 12'sd1574, 13'sd-2503}},
{{12'sd1562, 12'sd1586, 11'sd-565}, {12'sd1816, 11'sd-940, 8'sd93}, {13'sd2653, 12'sd1092, 13'sd-3628}},
{{13'sd-2290, 11'sd654, 11'sd-687}, {11'sd-552, 9'sd244, 12'sd1470}, {8'sd-115, 12'sd-1521, 10'sd-400}},
{{10'sd-472, 10'sd-453, 7'sd-52}, {13'sd3531, 12'sd-1654, 2'sd-1}, {12'sd1818, 11'sd-982, 13'sd3473}},
{{12'sd1650, 12'sd-1385, 11'sd-982}, {13'sd2171, 12'sd1222, 12'sd1250}, {12'sd-1397, 12'sd-2017, 13'sd2379}},
{{10'sd-317, 12'sd1968, 11'sd-750}, {9'sd-235, 11'sd882, 12'sd1208}, {12'sd-1112, 11'sd-524, 9'sd-171}},
{{13'sd2260, 6'sd20, 12'sd1746}, {13'sd2365, 13'sd-2214, 12'sd-1143}, {12'sd1597, 13'sd-2142, 11'sd808}},
{{13'sd2655, 10'sd355, 10'sd474}, {11'sd-886, 12'sd1591, 10'sd508}, {12'sd-1937, 13'sd-2798, 11'sd-838}},
{{12'sd1952, 13'sd2070, 10'sd426}, {12'sd-1852, 12'sd1564, 9'sd212}, {12'sd-1997, 12'sd-1377, 11'sd-821}},
{{12'sd1525, 12'sd1997, 12'sd1888}, {13'sd-2828, 12'sd1298, 12'sd-1866}, {12'sd1645, 9'sd160, 13'sd2613}},
{{7'sd-53, 10'sd-301, 12'sd1757}, {13'sd2663, 13'sd2088, 11'sd-847}, {11'sd-995, 11'sd-954, 13'sd4002}},
{{11'sd-543, 12'sd-1957, 13'sd-2163}, {13'sd-2168, 13'sd-2140, 12'sd1314}, {13'sd2298, 12'sd-1049, 11'sd-1003}},
{{13'sd2161, 12'sd1963, 10'sd427}, {13'sd2480, 12'sd1277, 12'sd-1751}, {11'sd-942, 13'sd2305, 7'sd33}},
{{8'sd111, 13'sd-2237, 10'sd335}, {12'sd1440, 10'sd456, 11'sd-957}, {13'sd-2197, 13'sd-2527, 12'sd1842}},
{{11'sd615, 12'sd1275, 12'sd1886}, {13'sd-3582, 12'sd1943, 11'sd-689}, {12'sd-2023, 13'sd-3016, 12'sd1293}},
{{12'sd1472, 12'sd1039, 13'sd2093}, {12'sd-1039, 12'sd1429, 13'sd2057}, {11'sd644, 12'sd1887, 12'sd1805}},
{{13'sd2789, 13'sd2571, 11'sd-755}, {13'sd2260, 12'sd-1070, 12'sd-1320}, {12'sd1959, 13'sd2707, 12'sd-1853}},
{{10'sd-311, 13'sd-2382, 13'sd-2804}, {12'sd-1568, 13'sd2180, 9'sd197}, {12'sd-1843, 11'sd-844, 11'sd-910}},
{{12'sd1924, 12'sd-1620, 11'sd-953}, {10'sd-479, 6'sd23, 11'sd-947}, {12'sd-1753, 10'sd389, 11'sd542}},
{{12'sd-1663, 13'sd2302, 12'sd-1487}, {13'sd-2238, 13'sd2053, 12'sd1044}, {13'sd-2371, 11'sd-568, 13'sd2062}},
{{12'sd-1055, 12'sd-1575, 9'sd132}, {10'sd-386, 10'sd-361, 11'sd-862}, {12'sd1118, 13'sd2573, 12'sd-1174}},
{{13'sd2556, 10'sd-445, 12'sd2027}, {13'sd2299, 8'sd-76, 7'sd33}, {13'sd-2101, 9'sd-175, 12'sd1252}},
{{6'sd28, 12'sd1389, 11'sd732}, {12'sd-1123, 9'sd-199, 12'sd-1875}, {13'sd-2293, 12'sd-1699, 11'sd-639}},
{{12'sd-1501, 8'sd115, 13'sd-2464}, {12'sd-1328, 12'sd-1741, 12'sd1509}, {13'sd-2425, 11'sd-765, 12'sd1682}},
{{12'sd-1675, 10'sd302, 12'sd1853}, {12'sd1757, 12'sd-1694, 12'sd1475}, {12'sd1957, 7'sd-63, 10'sd-373}},
{{12'sd-1815, 11'sd689, 10'sd326}, {11'sd614, 13'sd-2295, 12'sd-2046}, {11'sd-921, 13'sd2213, 10'sd-435}},
{{13'sd2343, 11'sd994, 12'sd1813}, {13'sd2139, 10'sd-375, 13'sd3230}, {13'sd2272, 13'sd2143, 13'sd2522}},
{{13'sd2351, 12'sd-1231, 12'sd-1265}, {13'sd2426, 12'sd1244, 13'sd2366}, {12'sd1227, 13'sd2077, 12'sd-1605}},
{{12'sd-1564, 12'sd1644, 11'sd-566}, {11'sd-545, 12'sd-1281, 12'sd1779}, {13'sd2305, 12'sd-1406, 13'sd2707}},
{{11'sd781, 11'sd-574, 8'sd124}, {13'sd-2196, 13'sd-2096, 11'sd-776}, {13'sd-2170, 11'sd-531, 11'sd539}},
{{11'sd1008, 12'sd1543, 13'sd-3522}, {13'sd-2906, 13'sd-2877, 13'sd-3463}, {13'sd-3744, 12'sd-1334, 13'sd-3740}},
{{11'sd596, 12'sd-1359, 13'sd2770}, {11'sd912, 7'sd-60, 12'sd-1202}, {9'sd-149, 12'sd-1827, 13'sd2484}},
{{13'sd-2072, 13'sd2578, 12'sd-1762}, {11'sd-656, 12'sd1551, 12'sd-1118}, {9'sd-178, 10'sd362, 10'sd327}},
{{12'sd1184, 12'sd1395, 12'sd1969}, {13'sd-2577, 13'sd-2194, 9'sd210}, {11'sd700, 12'sd-1373, 11'sd635}},
{{11'sd998, 13'sd-2748, 11'sd-654}, {11'sd650, 12'sd1655, 13'sd-2634}, {11'sd812, 13'sd2325, 8'sd91}},
{{10'sd-346, 11'sd761, 11'sd-740}, {12'sd1706, 12'sd1429, 11'sd828}, {10'sd-339, 13'sd2756, 12'sd-1182}},
{{13'sd3186, 10'sd-366, 11'sd800}, {13'sd3162, 13'sd3060, 12'sd1876}, {13'sd3808, 13'sd2061, 13'sd2339}},
{{12'sd1517, 12'sd-1758, 12'sd-1927}, {12'sd2017, 7'sd42, 10'sd449}, {11'sd820, 12'sd1772, 13'sd-2423}},
{{9'sd-211, 13'sd-2050, 11'sd848}, {13'sd-2117, 12'sd1437, 12'sd1446}, {11'sd-850, 13'sd-2423, 12'sd-1356}},
{{5'sd13, 9'sd253, 11'sd-690}, {12'sd1410, 12'sd-1066, 12'sd1608}, {12'sd-1934, 12'sd1721, 11'sd544}},
{{12'sd-1965, 8'sd103, 12'sd1374}, {12'sd-1964, 11'sd924, 12'sd-1188}, {12'sd-1555, 11'sd573, 11'sd851}},
{{13'sd2419, 13'sd-2547, 7'sd63}, {13'sd-2377, 12'sd-1855, 9'sd144}, {13'sd-2711, 10'sd288, 10'sd259}},
{{9'sd230, 10'sd286, 12'sd1085}, {9'sd161, 12'sd1741, 13'sd2726}, {13'sd-2422, 12'sd-1776, 13'sd-2546}},
{{13'sd-2783, 8'sd97, 12'sd1569}, {12'sd-1315, 13'sd2671, 12'sd1804}, {12'sd-1727, 13'sd-2605, 13'sd2424}},
{{13'sd-2305, 12'sd-1506, 7'sd-54}, {13'sd2356, 13'sd2308, 12'sd1490}, {9'sd209, 6'sd24, 12'sd1523}},
{{13'sd-3771, 13'sd-2725, 12'sd-1336}, {14'sd-4211, 11'sd903, 12'sd-1753}, {14'sd-4914, 12'sd-1049, 13'sd2517}},
{{13'sd2612, 12'sd1313, 13'sd-2220}, {13'sd-2531, 10'sd373, 11'sd-769}, {11'sd732, 11'sd-657, 10'sd-306}},
{{12'sd1049, 12'sd1582, 8'sd111}, {13'sd-2593, 12'sd1159, 13'sd-2597}, {11'sd977, 8'sd71, 12'sd1681}},
{{9'sd-169, 10'sd-355, 13'sd-2219}, {10'sd510, 13'sd-2209, 8'sd126}, {11'sd-522, 12'sd1113, 12'sd1028}},
{{13'sd-2305, 12'sd1673, 7'sd47}, {11'sd-730, 11'sd-752, 12'sd1397}, {13'sd-2652, 12'sd1810, 13'sd2194}},
{{13'sd3407, 9'sd-230, 13'sd2224}, {12'sd-1152, 12'sd-1157, 12'sd1294}, {13'sd3869, 13'sd2692, 10'sd-344}},
{{11'sd643, 12'sd1886, 12'sd-1759}, {13'sd2548, 13'sd2853, 10'sd-273}, {14'sd4718, 13'sd2299, 13'sd-3714}},
{{12'sd-1160, 11'sd577, 13'sd-2109}, {13'sd-3026, 9'sd-153, 10'sd296}, {11'sd-990, 13'sd2108, 12'sd-1773}},
{{13'sd2767, 10'sd503, 9'sd213}, {10'sd352, 10'sd310, 11'sd-843}, {10'sd-285, 12'sd1024, 13'sd-2232}},
{{13'sd-2679, 12'sd-1663, 11'sd804}, {12'sd-1410, 11'sd-877, 13'sd-2666}, {10'sd-308, 11'sd905, 9'sd254}},
{{12'sd-1442, 13'sd-2545, 10'sd-382}, {13'sd-2413, 9'sd194, 13'sd2381}, {13'sd2240, 13'sd-2506, 13'sd2488}},
{{13'sd-2894, 12'sd-1484, 13'sd2700}, {12'sd1785, 12'sd-1758, 9'sd-175}, {13'sd-3420, 12'sd1507, 11'sd737}}},
{
{{11'sd-945, 12'sd-1564, 12'sd1896}, {13'sd2245, 11'sd742, 13'sd3755}, {12'sd-1720, 12'sd1163, 10'sd-399}},
{{7'sd-38, 10'sd381, 12'sd-1604}, {12'sd1498, 12'sd-1700, 13'sd-2668}, {8'sd73, 12'sd1425, 13'sd-3284}},
{{12'sd1720, 10'sd377, 12'sd1730}, {9'sd-250, 11'sd-827, 13'sd-2226}, {12'sd-1581, 13'sd-2482, 12'sd1297}},
{{12'sd1610, 13'sd-2983, 12'sd-1395}, {10'sd-356, 13'sd2387, 11'sd851}, {10'sd508, 11'sd-947, 12'sd-1906}},
{{13'sd-3927, 6'sd-27, 12'sd1400}, {13'sd2239, 13'sd-2611, 12'sd-1285}, {13'sd3171, 10'sd499, 12'sd-1217}},
{{12'sd-1578, 13'sd2713, 11'sd-956}, {12'sd-1562, 12'sd1151, 11'sd-695}, {10'sd394, 11'sd601, 12'sd-1360}},
{{11'sd-715, 10'sd-387, 12'sd1647}, {12'sd1805, 11'sd567, 9'sd-220}, {12'sd1695, 9'sd176, 13'sd2613}},
{{13'sd-2690, 11'sd-986, 11'sd-514}, {14'sd-4294, 13'sd-2230, 13'sd-3590}, {11'sd599, 12'sd-1170, 11'sd-868}},
{{12'sd-1841, 12'sd-1886, 13'sd-2934}, {11'sd627, 13'sd-2495, 11'sd-916}, {9'sd-245, 9'sd193, 13'sd-2184}},
{{13'sd2263, 13'sd-2379, 13'sd2151}, {9'sd150, 11'sd731, 13'sd2810}, {10'sd-405, 13'sd2729, 12'sd-1790}},
{{12'sd1917, 13'sd3911, 14'sd4944}, {10'sd-378, 12'sd1469, 12'sd2047}, {13'sd2514, 13'sd-2121, 12'sd1130}},
{{12'sd-1212, 11'sd612, 12'sd1714}, {7'sd-56, 10'sd-416, 8'sd-97}, {13'sd-2281, 11'sd-881, 13'sd2729}},
{{11'sd542, 11'sd-721, 13'sd-2613}, {12'sd-2047, 12'sd-1524, 13'sd-3249}, {12'sd2013, 12'sd1078, 12'sd-1521}},
{{13'sd2532, 12'sd1430, 13'sd-2690}, {12'sd-1127, 12'sd-1372, 12'sd-2031}, {5'sd-11, 12'sd-1625, 13'sd-2632}},
{{12'sd1262, 12'sd1057, 11'sd580}, {12'sd-1973, 12'sd-1540, 12'sd1879}, {12'sd-1401, 11'sd-915, 10'sd-307}},
{{8'sd-127, 11'sd-993, 10'sd402}, {12'sd1702, 11'sd606, 11'sd-620}, {12'sd-1407, 13'sd3745, 9'sd-246}},
{{13'sd2676, 12'sd1750, 12'sd1158}, {10'sd-475, 12'sd1813, 12'sd-1065}, {13'sd3929, 14'sd4151, 13'sd2883}},
{{12'sd1114, 13'sd2815, 13'sd2329}, {13'sd-2425, 11'sd748, 6'sd-26}, {13'sd-3292, 12'sd1089, 11'sd747}},
{{13'sd-2956, 12'sd-1718, 13'sd-3515}, {10'sd-264, 13'sd-2423, 12'sd-1078}, {11'sd-774, 13'sd2412, 10'sd-337}},
{{11'sd-765, 13'sd-3194, 11'sd-640}, {11'sd-566, 13'sd-3784, 12'sd1446}, {11'sd912, 13'sd3877, 13'sd2996}},
{{4'sd4, 13'sd2559, 11'sd-585}, {10'sd-479, 12'sd1079, 10'sd-483}, {13'sd-2772, 13'sd-2817, 13'sd-3065}},
{{13'sd3179, 10'sd401, 11'sd522}, {13'sd2123, 9'sd145, 9'sd204}, {13'sd2773, 9'sd189, 12'sd1484}},
{{13'sd2241, 13'sd2218, 11'sd-984}, {12'sd-1558, 11'sd-753, 11'sd819}, {8'sd-82, 10'sd-391, 13'sd2673}},
{{13'sd-3242, 12'sd-1070, 12'sd1667}, {9'sd-252, 13'sd2438, 9'sd-243}, {11'sd-643, 13'sd2466, 10'sd321}},
{{12'sd1118, 12'sd-1044, 13'sd-2697}, {13'sd3260, 13'sd2283, 13'sd-2554}, {12'sd-1899, 11'sd-979, 13'sd-2298}},
{{12'sd-1435, 8'sd117, 13'sd-2094}, {12'sd1957, 13'sd-2863, 13'sd-2373}, {10'sd-496, 12'sd-1736, 12'sd1734}},
{{12'sd-1954, 11'sd-891, 12'sd1625}, {12'sd-1960, 13'sd2334, 12'sd-1686}, {10'sd-336, 11'sd-704, 9'sd182}},
{{13'sd-2641, 10'sd-275, 10'sd-329}, {11'sd-620, 11'sd-583, 13'sd-2482}, {13'sd-2278, 13'sd-2414, 12'sd1425}},
{{13'sd2428, 10'sd460, 11'sd580}, {12'sd-1362, 10'sd309, 11'sd-951}, {13'sd4074, 12'sd1933, 11'sd1007}},
{{12'sd1441, 9'sd195, 11'sd941}, {13'sd3820, 10'sd256, 12'sd1797}, {12'sd1165, 12'sd-1418, 13'sd2636}},
{{12'sd1797, 12'sd-2021, 12'sd-1641}, {11'sd-793, 12'sd-1253, 13'sd2208}, {10'sd-256, 12'sd1845, 13'sd2209}},
{{11'sd981, 13'sd-2087, 12'sd1524}, {10'sd265, 12'sd-1952, 13'sd-2166}, {11'sd820, 12'sd1811, 12'sd1919}},
{{12'sd-1981, 13'sd2392, 11'sd930}, {11'sd722, 11'sd719, 12'sd1162}, {11'sd-831, 10'sd-467, 13'sd2985}},
{{13'sd2487, 13'sd-2624, 10'sd-297}, {12'sd-1340, 13'sd-2159, 11'sd-851}, {12'sd1451, 10'sd369, 13'sd-2491}},
{{13'sd-2120, 13'sd-2968, 11'sd1016}, {10'sd470, 12'sd1335, 13'sd2725}, {12'sd-1332, 10'sd490, 12'sd1300}},
{{13'sd-2309, 12'sd1108, 11'sd736}, {13'sd2747, 13'sd2192, 7'sd44}, {11'sd981, 11'sd-597, 13'sd-3010}},
{{12'sd1613, 12'sd1227, 9'sd244}, {9'sd135, 11'sd904, 12'sd-1302}, {12'sd-2033, 13'sd-2594, 10'sd-415}},
{{10'sd463, 13'sd-2341, 13'sd2287}, {13'sd-2530, 9'sd186, 10'sd-371}, {11'sd-983, 12'sd1969, 12'sd1529}},
{{13'sd-3177, 12'sd-1985, 11'sd648}, {13'sd-2305, 13'sd-3283, 11'sd-948}, {11'sd-910, 13'sd-2652, 12'sd1801}},
{{10'sd-263, 11'sd639, 12'sd1853}, {12'sd-1169, 9'sd233, 13'sd2098}, {12'sd-1339, 11'sd776, 13'sd2650}},
{{13'sd2512, 13'sd2052, 11'sd-605}, {12'sd1862, 12'sd-1257, 11'sd856}, {13'sd2108, 10'sd333, 11'sd-939}},
{{13'sd-2858, 11'sd524, 12'sd1324}, {12'sd1660, 10'sd344, 13'sd2420}, {12'sd1511, 13'sd-2376, 12'sd1420}},
{{12'sd1727, 12'sd-1281, 10'sd-436}, {10'sd-381, 12'sd1931, 12'sd1414}, {13'sd2363, 10'sd-508, 12'sd-1071}},
{{12'sd1674, 12'sd1393, 12'sd1438}, {13'sd3687, 12'sd-1832, 12'sd-1270}, {11'sd-783, 12'sd-1859, 13'sd-3592}},
{{12'sd1566, 12'sd-1365, 10'sd324}, {12'sd1752, 13'sd2516, 10'sd476}, {13'sd2540, 10'sd-366, 12'sd1834}},
{{12'sd1533, 12'sd-1162, 13'sd-2528}, {13'sd-2799, 12'sd-2020, 12'sd-1028}, {10'sd443, 13'sd-3457, 12'sd1738}},
{{9'sd162, 13'sd3390, 12'sd-1215}, {11'sd737, 12'sd1901, 12'sd1027}, {13'sd2971, 13'sd2425, 12'sd1602}},
{{13'sd2674, 13'sd2845, 12'sd-1365}, {11'sd-826, 13'sd-2798, 11'sd-954}, {12'sd1228, 12'sd-1811, 11'sd679}},
{{9'sd161, 10'sd-404, 13'sd-2069}, {11'sd875, 11'sd777, 10'sd374}, {13'sd-2132, 13'sd2148, 11'sd874}},
{{10'sd-379, 11'sd-589, 12'sd1168}, {11'sd850, 11'sd-761, 12'sd-1146}, {12'sd1071, 11'sd-608, 12'sd1210}},
{{12'sd1904, 13'sd-2454, 12'sd-1468}, {13'sd2671, 12'sd-1998, 9'sd-235}, {12'sd1619, 13'sd2858, 10'sd-396}},
{{12'sd-1235, 13'sd-2349, 13'sd2254}, {13'sd-2151, 12'sd1684, 12'sd-1249}, {5'sd12, 12'sd1848, 11'sd1012}},
{{11'sd908, 12'sd1844, 13'sd3210}, {8'sd86, 12'sd1120, 11'sd681}, {12'sd-1775, 12'sd-1704, 12'sd-1930}},
{{13'sd2179, 12'sd1623, 13'sd-2078}, {12'sd-1934, 12'sd-1269, 10'sd-427}, {12'sd-1878, 11'sd-833, 12'sd1563}},
{{11'sd-532, 13'sd-2071, 13'sd2755}, {12'sd1124, 12'sd-1058, 13'sd2309}, {11'sd777, 13'sd2523, 10'sd-425}},
{{12'sd-1620, 13'sd-2255, 12'sd1416}, {12'sd1379, 9'sd201, 11'sd-962}, {12'sd-2026, 12'sd-1422, 12'sd-1089}},
{{12'sd1712, 11'sd-970, 13'sd-2270}, {11'sd823, 12'sd-1080, 13'sd-3022}, {10'sd-444, 12'sd2033, 10'sd-379}},
{{10'sd372, 10'sd-387, 12'sd1855}, {13'sd-2473, 12'sd1113, 11'sd602}, {12'sd-1283, 13'sd-2107, 11'sd943}},
{{13'sd2403, 11'sd1023, 13'sd3373}, {10'sd309, 13'sd3577, 14'sd5160}, {13'sd-3897, 10'sd463, 13'sd2640}},
{{11'sd-669, 12'sd-1903, 13'sd-2255}, {13'sd2086, 12'sd1661, 12'sd1921}, {12'sd1535, 11'sd798, 12'sd1138}},
{{11'sd536, 13'sd-2380, 13'sd2065}, {11'sd882, 9'sd152, 12'sd1844}, {13'sd-2412, 9'sd178, 12'sd1705}},
{{9'sd248, 12'sd-1277, 10'sd317}, {13'sd3314, 10'sd501, 9'sd229}, {13'sd2225, 11'sd-718, 13'sd2468}},
{{12'sd-1388, 12'sd-1697, 10'sd-339}, {13'sd2986, 12'sd1741, 10'sd-453}, {12'sd-2000, 12'sd-1583, 12'sd-1946}},
{{13'sd-2732, 12'sd1940, 13'sd3811}, {12'sd-1409, 12'sd-1947, 13'sd2891}, {13'sd2461, 13'sd2547, 12'sd-1036}}},
{
{{11'sd793, 12'sd-1568, 12'sd1185}, {12'sd-1178, 9'sd215, 12'sd1843}, {12'sd-1650, 11'sd656, 10'sd431}},
{{13'sd-2941, 13'sd-2836, 12'sd-1688}, {13'sd-2424, 11'sd552, 11'sd-699}, {13'sd2091, 12'sd1408, 12'sd1290}},
{{12'sd-1115, 12'sd-1222, 11'sd764}, {12'sd-1992, 12'sd-1211, 12'sd-1367}, {11'sd828, 11'sd-709, 10'sd-510}},
{{13'sd-2204, 13'sd2135, 13'sd2391}, {11'sd-576, 11'sd-917, 13'sd2279}, {12'sd-1357, 13'sd2841, 13'sd-2194}},
{{10'sd267, 12'sd-1894, 12'sd-1689}, {13'sd2185, 11'sd882, 12'sd-1867}, {11'sd620, 13'sd-2586, 13'sd-3187}},
{{12'sd1038, 13'sd-2420, 13'sd2687}, {8'sd76, 11'sd-618, 13'sd2460}, {13'sd2231, 11'sd973, 13'sd2350}},
{{10'sd299, 12'sd1732, 12'sd1099}, {12'sd-1316, 13'sd-2345, 11'sd638}, {9'sd-181, 13'sd2233, 10'sd458}},
{{11'sd-574, 12'sd1192, 11'sd-1023}, {13'sd2564, 12'sd1887, 9'sd204}, {12'sd1603, 10'sd295, 13'sd2160}},
{{12'sd-1334, 13'sd-2407, 12'sd1044}, {11'sd717, 12'sd1315, 12'sd1665}, {12'sd1772, 10'sd-401, 12'sd1339}},
{{12'sd-1744, 11'sd537, 13'sd2748}, {9'sd-210, 10'sd-510, 13'sd-3049}, {13'sd2373, 11'sd606, 12'sd1966}},
{{13'sd3993, 12'sd-1233, 12'sd-1236}, {13'sd3681, 13'sd2148, 12'sd1557}, {13'sd2381, 11'sd814, 10'sd481}},
{{11'sd528, 13'sd2272, 11'sd-604}, {13'sd2337, 12'sd1857, 9'sd237}, {13'sd-3150, 13'sd2204, 13'sd-3072}},
{{12'sd-1942, 13'sd-2290, 11'sd700}, {12'sd-1567, 13'sd-2585, 13'sd2235}, {13'sd2101, 13'sd2483, 12'sd-1976}},
{{11'sd648, 10'sd-413, 9'sd159}, {13'sd2665, 12'sd-1956, 10'sd458}, {8'sd102, 11'sd-732, 8'sd88}},
{{13'sd-2593, 12'sd-1567, 13'sd2139}, {12'sd-1367, 11'sd520, 12'sd1478}, {12'sd-1819, 11'sd747, 12'sd1636}},
{{12'sd2027, 11'sd-668, 12'sd1037}, {9'sd192, 12'sd-1041, 11'sd-609}, {10'sd328, 11'sd675, 8'sd-111}},
{{12'sd1622, 12'sd-2040, 9'sd173}, {7'sd-57, 11'sd-804, 12'sd-1332}, {12'sd-1433, 8'sd66, 12'sd-1665}},
{{13'sd-2102, 13'sd-3078, 11'sd-643}, {12'sd-1730, 13'sd-2414, 12'sd-1590}, {13'sd-2134, 11'sd-574, 10'sd-405}},
{{12'sd-1817, 13'sd2765, 11'sd-590}, {10'sd415, 13'sd3048, 12'sd1170}, {13'sd-2632, 12'sd1553, 12'sd-1381}},
{{13'sd2342, 12'sd-1497, 12'sd-1087}, {12'sd-1198, 10'sd-391, 10'sd-429}, {13'sd4012, 13'sd2061, 11'sd674}},
{{12'sd1210, 12'sd-1554, 8'sd-99}, {13'sd-2501, 12'sd-1252, 12'sd1445}, {12'sd-1342, 12'sd-1122, 12'sd2031}},
{{14'sd-4955, 12'sd-1445, 12'sd-1559}, {12'sd-1215, 13'sd-2675, 13'sd2166}, {11'sd984, 11'sd892, 13'sd2333}},
{{12'sd1666, 11'sd574, 12'sd1898}, {12'sd-1280, 13'sd-2350, 13'sd2333}, {11'sd-612, 11'sd780, 11'sd963}},
{{11'sd-962, 12'sd-2046, 10'sd451}, {12'sd2044, 10'sd368, 12'sd-1653}, {10'sd349, 11'sd-750, 11'sd864}},
{{11'sd825, 12'sd1647, 12'sd-1204}, {13'sd-2402, 11'sd-552, 12'sd1682}, {14'sd-5459, 13'sd-3880, 12'sd-1175}},
{{12'sd1827, 13'sd2475, 11'sd-622}, {10'sd486, 13'sd2478, 12'sd-1135}, {12'sd-1919, 13'sd-2207, 12'sd-1991}},
{{12'sd1039, 13'sd-2474, 13'sd-2127}, {12'sd-1621, 10'sd296, 10'sd-307}, {12'sd-1596, 11'sd-704, 11'sd818}},
{{12'sd1341, 13'sd2404, 10'sd437}, {13'sd-2202, 12'sd1922, 12'sd1398}, {13'sd2664, 12'sd-1370, 7'sd-34}},
{{12'sd-1459, 13'sd-2987, 10'sd-280}, {11'sd718, 12'sd-1033, 12'sd-1883}, {13'sd2873, 12'sd1649, 10'sd-260}},
{{13'sd-2230, 12'sd-1222, 9'sd-241}, {12'sd1663, 12'sd1344, 12'sd-1173}, {5'sd14, 13'sd2493, 10'sd269}},
{{12'sd-1505, 12'sd1439, 12'sd1994}, {10'sd-435, 12'sd1279, 12'sd1788}, {12'sd-1357, 12'sd-1945, 11'sd806}},
{{12'sd1776, 9'sd-199, 13'sd2230}, {12'sd-1714, 12'sd1441, 13'sd-2566}, {10'sd-275, 13'sd-2900, 10'sd-457}},
{{10'sd-489, 11'sd720, 11'sd768}, {12'sd1400, 12'sd-1872, 13'sd-2140}, {12'sd1469, 11'sd-644, 12'sd1978}},
{{12'sd1872, 13'sd-2813, 13'sd-2372}, {13'sd-2360, 12'sd1567, 11'sd-681}, {12'sd1106, 12'sd1396, 12'sd1765}},
{{13'sd2787, 10'sd408, 12'sd1843}, {12'sd1294, 13'sd-2061, 11'sd820}, {13'sd-2099, 12'sd-1098, 10'sd342}},
{{11'sd-942, 12'sd1330, 13'sd-2070}, {13'sd2052, 9'sd-129, 10'sd-348}, {13'sd-2555, 9'sd191, 13'sd-2175}},
{{13'sd-3186, 13'sd-3322, 10'sd-300}, {11'sd-846, 12'sd-1985, 12'sd1110}, {13'sd2157, 13'sd2093, 12'sd-1524}},
{{13'sd3205, 12'sd1100, 12'sd-1384}, {8'sd83, 12'sd-1260, 13'sd3089}, {11'sd731, 14'sd-4098, 14'sd-4376}},
{{13'sd3135, 13'sd2683, 13'sd2923}, {13'sd2843, 12'sd1731, 10'sd319}, {12'sd-2021, 12'sd1281, 13'sd-2123}},
{{12'sd1798, 12'sd-1531, 11'sd-827}, {11'sd985, 11'sd-562, 11'sd-624}, {13'sd-2521, 13'sd-2670, 9'sd-142}},
{{13'sd-2464, 13'sd2668, 12'sd1567}, {12'sd1438, 11'sd-911, 12'sd-1424}, {12'sd1639, 13'sd-3023, 12'sd1645}},
{{12'sd-1476, 13'sd2538, 12'sd1072}, {11'sd-598, 13'sd2843, 13'sd2633}, {12'sd1119, 8'sd77, 12'sd-1788}},
{{9'sd-135, 10'sd-289, 13'sd2760}, {13'sd-2411, 9'sd-150, 6'sd-19}, {11'sd950, 13'sd2953, 13'sd2622}},
{{10'sd-507, 12'sd1673, 11'sd-589}, {7'sd52, 13'sd2640, 12'sd-1440}, {13'sd-3364, 13'sd2177, 12'sd-1983}},
{{12'sd-1242, 9'sd-166, 11'sd-806}, {12'sd-1537, 11'sd987, 10'sd-448}, {13'sd2659, 11'sd971, 10'sd334}},
{{13'sd-3383, 13'sd-2664, 12'sd-1479}, {11'sd633, 8'sd-98, 12'sd1030}, {13'sd2609, 12'sd1482, 11'sd-707}},
{{12'sd1976, 12'sd1662, 12'sd1059}, {12'sd-1625, 12'sd1825, 11'sd-548}, {13'sd-2727, 12'sd-1824, 12'sd-1612}},
{{12'sd-1644, 12'sd-1267, 12'sd1535}, {9'sd-139, 12'sd-1809, 11'sd592}, {10'sd-356, 6'sd23, 11'sd712}},
{{12'sd1466, 12'sd1573, 10'sd499}, {12'sd-1334, 12'sd-1355, 13'sd-2702}, {13'sd-2911, 13'sd2390, 12'sd1115}},
{{10'sd263, 12'sd-1833, 12'sd-1139}, {12'sd-1067, 6'sd-22, 12'sd-1841}, {9'sd-252, 12'sd1528, 9'sd220}},
{{13'sd2050, 11'sd625, 7'sd59}, {12'sd-1786, 12'sd2030, 12'sd-1442}, {10'sd317, 12'sd1094, 13'sd-2426}},
{{12'sd1192, 13'sd2723, 12'sd-1580}, {11'sd680, 11'sd554, 12'sd1162}, {13'sd-2387, 12'sd-1381, 12'sd1831}},
{{13'sd-2648, 11'sd-514, 13'sd-2277}, {13'sd-3791, 12'sd1646, 13'sd2235}, {9'sd140, 12'sd-1184, 13'sd2187}},
{{11'sd1009, 12'sd1109, 12'sd-1271}, {13'sd2084, 10'sd-308, 10'sd-365}, {11'sd782, 10'sd-336, 12'sd-1326}},
{{9'sd254, 10'sd374, 13'sd2179}, {11'sd818, 12'sd1669, 12'sd1904}, {12'sd1606, 13'sd-2939, 12'sd-2034}},
{{10'sd422, 11'sd-610, 11'sd694}, {8'sd-103, 13'sd-2221, 13'sd-2559}, {13'sd3134, 13'sd2236, 13'sd2396}},
{{12'sd1717, 13'sd-3148, 9'sd135}, {13'sd2409, 12'sd-1707, 13'sd2970}, {12'sd1685, 12'sd-1824, 13'sd2355}},
{{12'sd1243, 13'sd2348, 10'sd-332}, {11'sd-797, 13'sd2193, 11'sd-898}, {12'sd-1873, 11'sd903, 12'sd1458}},
{{13'sd2675, 13'sd-4002, 12'sd-1892}, {13'sd2526, 12'sd-1558, 10'sd303}, {13'sd3562, 13'sd2350, 10'sd-380}},
{{12'sd1655, 12'sd-1565, 12'sd-1917}, {8'sd-94, 13'sd2600, 12'sd1694}, {11'sd1002, 7'sd-59, 13'sd2491}},
{{12'sd1705, 11'sd552, 11'sd-690}, {11'sd516, 13'sd-2270, 12'sd-1671}, {13'sd-2357, 12'sd-1562, 10'sd429}},
{{12'sd1956, 10'sd313, 10'sd418}, {10'sd-265, 12'sd-1727, 12'sd1407}, {7'sd-34, 13'sd2227, 13'sd-2669}},
{{10'sd411, 12'sd1462, 12'sd1531}, {12'sd1575, 12'sd2045, 11'sd-965}, {13'sd-2069, 13'sd-2358, 12'sd1179}},
{{9'sd134, 13'sd2259, 10'sd309}, {12'sd1619, 13'sd-2143, 12'sd-1047}, {13'sd-3282, 12'sd1550, 11'sd626}}},
{
{{13'sd-2081, 10'sd384, 11'sd805}, {12'sd-1406, 12'sd-1294, 14'sd4281}, {10'sd395, 10'sd360, 13'sd3286}},
{{13'sd-2470, 12'sd-1518, 11'sd-773}, {10'sd410, 12'sd1644, 13'sd2149}, {13'sd2954, 11'sd-1004, 11'sd-610}},
{{14'sd4252, 9'sd168, 12'sd1086}, {13'sd3325, 12'sd-1365, 9'sd174}, {8'sd68, 12'sd-1723, 13'sd-2475}},
{{13'sd-2991, 12'sd-2008, 12'sd1236}, {12'sd-1376, 11'sd761, 12'sd1863}, {11'sd-1016, 12'sd-1518, 12'sd1186}},
{{13'sd-3522, 13'sd2225, 13'sd-2114}, {8'sd-70, 13'sd2644, 12'sd-1304}, {12'sd1887, 12'sd-1236, 11'sd863}},
{{10'sd-272, 12'sd-1040, 11'sd-630}, {13'sd2313, 12'sd2006, 12'sd1405}, {12'sd-1889, 5'sd11, 11'sd-728}},
{{12'sd-1247, 12'sd-1519, 12'sd1129}, {14'sd-4139, 11'sd-814, 12'sd-1256}, {9'sd249, 11'sd-884, 1'sd0}},
{{13'sd-2095, 14'sd-4457, 12'sd1854}, {10'sd265, 14'sd-4128, 12'sd1230}, {12'sd1767, 11'sd-614, 13'sd3770}},
{{10'sd-317, 8'sd-66, 14'sd4528}, {11'sd-699, 12'sd1578, 10'sd385}, {12'sd-1924, 9'sd-220, 11'sd-1023}},
{{13'sd2703, 5'sd-14, 13'sd-2093}, {11'sd-1022, 11'sd-1003, 12'sd-1882}, {11'sd862, 11'sd685, 13'sd2104}},
{{11'sd718, 14'sd4998, 11'sd678}, {12'sd1683, 14'sd5398, 9'sd201}, {13'sd2877, 12'sd1535, 8'sd-96}},
{{11'sd-971, 7'sd-62, 13'sd-2517}, {13'sd-2639, 10'sd367, 13'sd3001}, {12'sd-1859, 12'sd1797, 13'sd2591}},
{{11'sd-535, 13'sd-2561, 13'sd-2775}, {8'sd118, 13'sd-2678, 12'sd-1375}, {5'sd-9, 12'sd-1064, 12'sd-1097}},
{{9'sd-220, 9'sd-243, 10'sd-467}, {11'sd-882, 13'sd2447, 12'sd-1841}, {12'sd-1527, 13'sd3002, 13'sd3830}},
{{7'sd44, 12'sd1782, 11'sd534}, {11'sd720, 13'sd2461, 11'sd581}, {12'sd-1508, 10'sd489, 11'sd943}},
{{12'sd-1688, 12'sd1139, 13'sd-3467}, {13'sd-3015, 13'sd-3244, 13'sd-2170}, {11'sd567, 7'sd36, 13'sd3284}},
{{11'sd-606, 12'sd-1834, 13'sd-2971}, {11'sd942, 12'sd-1707, 8'sd82}, {12'sd1650, 12'sd1398, 7'sd-63}},
{{13'sd3056, 13'sd2272, 12'sd1389}, {12'sd1400, 13'sd2235, 13'sd-2611}, {11'sd-851, 11'sd984, 14'sd-4598}},
{{13'sd-3852, 12'sd-1594, 10'sd418}, {11'sd-985, 12'sd-1704, 13'sd2048}, {9'sd170, 13'sd2424, 13'sd3036}},
{{12'sd-1602, 13'sd3464, 12'sd-1250}, {12'sd1658, 13'sd3439, 12'sd1579}, {11'sd566, 11'sd661, 11'sd598}},
{{9'sd168, 12'sd1325, 12'sd-1897}, {12'sd1520, 11'sd-717, 12'sd1937}, {9'sd-246, 12'sd-1388, 7'sd55}},
{{12'sd1667, 13'sd-3509, 12'sd-1625}, {14'sd4504, 10'sd505, 11'sd-802}, {14'sd5620, 12'sd1782, 10'sd406}},
{{13'sd3886, 11'sd-583, 12'sd-1929}, {13'sd2429, 13'sd-2266, 11'sd990}, {13'sd2930, 10'sd-382, 10'sd447}},
{{8'sd-101, 13'sd2065, 10'sd-303}, {9'sd-195, 11'sd-911, 12'sd1270}, {13'sd-2319, 13'sd-3142, 13'sd-3432}},
{{10'sd-275, 14'sd-4346, 13'sd-2744}, {13'sd2065, 12'sd-1622, 13'sd2600}, {10'sd276, 13'sd-3769, 11'sd-805}},
{{11'sd-970, 12'sd1986, 12'sd-1257}, {13'sd-2877, 11'sd-655, 10'sd492}, {12'sd-1106, 12'sd-2046, 13'sd3731}},
{{12'sd-1775, 11'sd979, 13'sd2217}, {13'sd-3241, 13'sd2164, 11'sd-1003}, {12'sd-1863, 6'sd-27, 10'sd-265}},
{{9'sd165, 11'sd968, 13'sd3027}, {10'sd440, 12'sd-1227, 11'sd-1004}, {13'sd2234, 11'sd564, 11'sd898}},
{{12'sd1712, 12'sd-1882, 12'sd-1105}, {13'sd-2941, 13'sd-2673, 13'sd-3265}, {13'sd3570, 12'sd1416, 13'sd-2494}},
{{12'sd1731, 10'sd299, 13'sd-3007}, {10'sd468, 12'sd-1322, 12'sd2023}, {13'sd2935, 12'sd-1702, 13'sd-2489}},
{{11'sd735, 10'sd-401, 12'sd-1138}, {11'sd659, 7'sd-35, 13'sd-2805}, {11'sd-776, 5'sd-14, 10'sd276}},
{{12'sd1522, 12'sd1115, 13'sd2196}, {12'sd-1809, 13'sd2517, 11'sd722}, {12'sd-1526, 12'sd1919, 14'sd4574}},
{{10'sd421, 9'sd180, 12'sd-1916}, {13'sd3776, 12'sd-1504, 13'sd-2760}, {11'sd819, 11'sd-818, 12'sd-1178}},
{{13'sd2561, 10'sd333, 12'sd1257}, {13'sd3323, 12'sd1325, 11'sd887}, {13'sd2375, 9'sd-160, 13'sd-3808}},
{{13'sd-3027, 11'sd-821, 13'sd-3299}, {10'sd-262, 13'sd3754, 10'sd-431}, {11'sd-764, 12'sd1677, 13'sd2326}},
{{13'sd-2582, 11'sd541, 12'sd1165}, {12'sd-1562, 11'sd-565, 10'sd292}, {13'sd2084, 11'sd-665, 11'sd-651}},
{{13'sd2878, 8'sd99, 11'sd728}, {12'sd1270, 9'sd-199, 13'sd-2467}, {11'sd802, 13'sd-2525, 9'sd-204}},
{{14'sd-4343, 12'sd1344, 11'sd-814}, {6'sd19, 12'sd2028, 10'sd469}, {9'sd-188, 10'sd390, 13'sd2792}},
{{13'sd-2238, 13'sd2820, 10'sd317}, {11'sd-537, 9'sd210, 11'sd-1013}, {12'sd1867, 10'sd298, 13'sd2242}},
{{13'sd-3280, 12'sd1074, 12'sd-1696}, {12'sd1770, 13'sd2155, 12'sd-1627}, {10'sd-335, 13'sd2778, 9'sd-247}},
{{12'sd-1855, 12'sd1141, 7'sd57}, {10'sd-439, 13'sd-2379, 12'sd1696}, {8'sd127, 12'sd-1648, 12'sd-1028}},
{{13'sd-3717, 11'sd-759, 11'sd-916}, {12'sd-1321, 7'sd53, 12'sd1942}, {12'sd2023, 12'sd-1129, 12'sd1330}},
{{10'sd337, 11'sd-550, 12'sd1251}, {11'sd868, 13'sd3360, 13'sd2482}, {11'sd-546, 11'sd698, 12'sd1407}},
{{10'sd-434, 11'sd-523, 13'sd2169}, {11'sd-866, 11'sd-950, 12'sd1727}, {11'sd-783, 10'sd405, 13'sd3217}},
{{10'sd327, 10'sd-435, 12'sd1240}, {12'sd1544, 13'sd2285, 11'sd-597}, {9'sd151, 12'sd-1668, 13'sd-3600}},
{{12'sd1086, 13'sd2127, 12'sd-1268}, {12'sd1949, 8'sd86, 11'sd-906}, {13'sd2304, 10'sd-371, 13'sd-3768}},
{{12'sd-1578, 12'sd1119, 11'sd723}, {11'sd-715, 13'sd-2249, 10'sd-344}, {13'sd2191, 12'sd-1584, 11'sd-877}},
{{12'sd1292, 11'sd857, 11'sd-695}, {13'sd3102, 13'sd2566, 12'sd2029}, {12'sd1149, 12'sd1081, 12'sd-2047}},
{{11'sd-597, 11'sd-768, 12'sd1644}, {12'sd1410, 12'sd-1411, 12'sd1360}, {11'sd768, 10'sd334, 7'sd38}},
{{12'sd1297, 13'sd-3097, 13'sd-2157}, {11'sd-986, 10'sd346, 12'sd-1044}, {6'sd26, 12'sd-1553, 10'sd-427}},
{{11'sd802, 9'sd-229, 13'sd2164}, {10'sd493, 11'sd-726, 13'sd2084}, {11'sd645, 11'sd-999, 12'sd-1116}},
{{11'sd656, 13'sd-2523, 12'sd-1902}, {13'sd2452, 12'sd2046, 12'sd1761}, {13'sd-2111, 12'sd1409, 13'sd-2586}},
{{6'sd20, 12'sd-1256, 11'sd934}, {12'sd1364, 12'sd-1074, 10'sd353}, {13'sd2899, 10'sd-342, 13'sd-3849}},
{{12'sd1836, 12'sd2041, 10'sd-263}, {11'sd-989, 13'sd2307, 11'sd925}, {10'sd-292, 11'sd-1001, 12'sd-1159}},
{{12'sd-1239, 13'sd-2079, 13'sd-2899}, {13'sd2246, 13'sd2148, 11'sd-985}, {10'sd-394, 11'sd626, 9'sd-253}},
{{12'sd1720, 12'sd-1662, 11'sd-755}, {9'sd-164, 8'sd-116, 12'sd-1026}, {11'sd-947, 13'sd-2753, 13'sd-3906}},
{{10'sd309, 12'sd1816, 13'sd-2587}, {8'sd-82, 10'sd-456, 12'sd1329}, {13'sd-2318, 12'sd-1722, 11'sd-748}},
{{12'sd-1445, 11'sd-793, 11'sd-991}, {14'sd-5002, 12'sd1494, 13'sd3045}, {14'sd-5735, 10'sd-450, 11'sd-618}},
{{13'sd2580, 12'sd1790, 13'sd3707}, {14'sd-4259, 5'sd8, 13'sd4025}, {13'sd-3146, 12'sd-1035, 14'sd6250}},
{{13'sd-3199, 11'sd556, 12'sd-1421}, {12'sd-1951, 12'sd1833, 13'sd2574}, {13'sd2836, 12'sd1489, 11'sd751}},
{{12'sd-1765, 13'sd-4049, 13'sd-2572}, {11'sd-868, 12'sd1167, 13'sd2405}, {12'sd1628, 13'sd2174, 11'sd-708}},
{{12'sd-1596, 13'sd-2501, 10'sd350}, {12'sd1046, 13'sd-2568, 11'sd-769}, {13'sd2622, 12'sd1472, 12'sd1691}},
{{12'sd-1124, 12'sd1973, 12'sd1971}, {11'sd-866, 11'sd-795, 10'sd-492}, {11'sd946, 12'sd2005, 13'sd3361}},
{{13'sd-2210, 11'sd958, 13'sd2315}, {13'sd2440, 10'sd347, 13'sd2432}, {12'sd-1792, 12'sd-2005, 12'sd-1585}}},
{
{{11'sd-952, 13'sd2204, 13'sd2263}, {12'sd1418, 12'sd1836, 12'sd1068}, {13'sd-2144, 13'sd3211, 13'sd2882}},
{{10'sd473, 13'sd2628, 10'sd-425}, {10'sd-271, 12'sd1389, 12'sd1997}, {12'sd-1975, 11'sd-635, 11'sd800}},
{{12'sd1076, 12'sd-1123, 13'sd-3366}, {13'sd-2290, 10'sd364, 12'sd-1854}, {12'sd1737, 9'sd189, 12'sd1856}},
{{11'sd892, 12'sd1230, 13'sd-2178}, {11'sd664, 13'sd2227, 8'sd-68}, {10'sd270, 12'sd1042, 10'sd-440}},
{{11'sd-740, 9'sd206, 12'sd1605}, {13'sd2641, 12'sd-1847, 12'sd1175}, {12'sd1518, 13'sd2573, 11'sd666}},
{{13'sd2304, 10'sd-294, 12'sd-1657}, {11'sd650, 8'sd-104, 13'sd-2304}, {8'sd76, 10'sd-448, 12'sd-1477}},
{{11'sd672, 11'sd832, 11'sd645}, {12'sd1548, 12'sd1880, 11'sd703}, {9'sd172, 11'sd786, 11'sd691}},
{{10'sd389, 12'sd1428, 13'sd-2110}, {12'sd1151, 12'sd-1212, 13'sd2085}, {13'sd-2656, 8'sd127, 10'sd-372}},
{{12'sd-1096, 12'sd-1471, 11'sd874}, {11'sd-806, 13'sd-2473, 11'sd526}, {12'sd1664, 13'sd-2936, 12'sd1644}},
{{13'sd2726, 11'sd-704, 12'sd2024}, {11'sd997, 11'sd-747, 12'sd1341}, {13'sd2288, 12'sd1764, 13'sd2661}},
{{14'sd-5115, 13'sd-3830, 11'sd939}, {12'sd-1571, 13'sd-3082, 12'sd1250}, {14'sd-4365, 11'sd-951, 12'sd-1923}},
{{10'sd276, 11'sd-791, 11'sd787}, {12'sd1163, 12'sd-1814, 10'sd-350}, {12'sd-1797, 13'sd-2154, 13'sd-2048}},
{{11'sd-524, 12'sd1102, 11'sd785}, {11'sd-588, 6'sd26, 12'sd1259}, {13'sd3403, 13'sd2766, 12'sd-1843}},
{{12'sd-1298, 13'sd-2797, 11'sd-603}, {12'sd2026, 13'sd-2738, 11'sd-924}, {8'sd102, 12'sd-1409, 13'sd-2262}},
{{12'sd-1217, 12'sd1106, 8'sd125}, {12'sd-1680, 13'sd-2723, 12'sd-1461}, {12'sd2018, 12'sd-1056, 10'sd-342}},
{{10'sd303, 11'sd-765, 13'sd2464}, {13'sd-2470, 10'sd-307, 7'sd-50}, {11'sd-988, 11'sd-736, 10'sd-470}},
{{12'sd1275, 11'sd-776, 12'sd2021}, {11'sd656, 13'sd-2064, 11'sd-932}, {13'sd3044, 12'sd-1142, 8'sd106}},
{{11'sd524, 13'sd3279, 12'sd-1647}, {10'sd-336, 11'sd-755, 8'sd-121}, {13'sd2907, 8'sd-67, 13'sd-3038}},
{{12'sd1410, 13'sd2114, 13'sd-2483}, {11'sd-668, 13'sd-2532, 13'sd2537}, {9'sd-157, 11'sd871, 11'sd-909}},
{{12'sd-1469, 13'sd-2196, 12'sd1362}, {12'sd1312, 13'sd-2399, 13'sd3040}, {10'sd343, 12'sd1709, 12'sd1932}},
{{13'sd-2129, 12'sd1272, 12'sd2030}, {12'sd1363, 13'sd2272, 12'sd1836}, {11'sd-991, 11'sd927, 13'sd-2389}},
{{12'sd1801, 13'sd-2504, 12'sd1590}, {10'sd-277, 12'sd1120, 13'sd-3108}, {10'sd460, 13'sd2362, 9'sd-208}},
{{10'sd348, 12'sd-1118, 12'sd1665}, {12'sd1450, 12'sd-1312, 10'sd418}, {12'sd1717, 13'sd2091, 13'sd2080}},
{{13'sd-3094, 11'sd-771, 13'sd2100}, {13'sd-2905, 12'sd-1212, 12'sd-1275}, {13'sd-3366, 12'sd1333, 13'sd-2122}},
{{11'sd548, 13'sd3935, 12'sd1680}, {10'sd-438, 11'sd1019, 12'sd1320}, {13'sd2292, 13'sd2743, 12'sd1944}},
{{11'sd-700, 12'sd1990, 12'sd1418}, {13'sd2693, 11'sd542, 10'sd477}, {9'sd-174, 12'sd1138, 9'sd231}},
{{12'sd-1797, 12'sd1557, 12'sd1267}, {13'sd2395, 12'sd2030, 12'sd-1337}, {13'sd-2560, 10'sd-305, 12'sd1038}},
{{11'sd-540, 13'sd-2076, 10'sd-481}, {13'sd2557, 12'sd-1140, 12'sd1046}, {11'sd-926, 9'sd193, 12'sd-1793}},
{{12'sd-1485, 12'sd1575, 10'sd281}, {12'sd-1696, 12'sd-1758, 13'sd-2508}, {12'sd-1220, 13'sd2402, 13'sd-2139}},
{{8'sd68, 12'sd-1527, 11'sd-736}, {12'sd1960, 13'sd-3043, 12'sd1513}, {13'sd2240, 12'sd-1090, 13'sd2131}},
{{12'sd-1406, 7'sd-44, 10'sd-392}, {12'sd-1817, 12'sd1872, 11'sd-817}, {8'sd74, 12'sd1747, 13'sd2556}},
{{12'sd-1512, 12'sd1248, 11'sd-591}, {12'sd1469, 9'sd220, 12'sd-1538}, {10'sd-290, 10'sd-447, 11'sd989}},
{{13'sd-2100, 12'sd-1639, 13'sd-2073}, {12'sd1523, 11'sd-754, 12'sd-1262}, {12'sd1414, 12'sd-2014, 11'sd-586}},
{{13'sd2723, 12'sd1345, 11'sd540}, {13'sd2482, 10'sd-382, 12'sd-1812}, {8'sd112, 12'sd1483, 6'sd-29}},
{{12'sd1393, 13'sd-2452, 10'sd411}, {13'sd-2317, 12'sd1569, 12'sd-1317}, {12'sd-2030, 12'sd-1304, 11'sd-735}},
{{12'sd1846, 11'sd823, 12'sd-1778}, {12'sd-1313, 12'sd-1317, 9'sd-164}, {13'sd-2465, 7'sd-43, 12'sd1852}},
{{13'sd2111, 12'sd-1964, 11'sd-912}, {11'sd822, 7'sd52, 11'sd-602}, {12'sd1831, 5'sd15, 12'sd-1682}},
{{13'sd-2960, 11'sd-886, 12'sd-1738}, {13'sd2321, 12'sd-1106, 12'sd1176}, {10'sd342, 12'sd1329, 13'sd2307}},
{{12'sd-1324, 12'sd1713, 12'sd1901}, {11'sd880, 12'sd-1840, 13'sd2508}, {13'sd2746, 12'sd1375, 13'sd2459}},
{{12'sd-1115, 12'sd1441, 11'sd792}, {10'sd439, 7'sd41, 10'sd316}, {12'sd1512, 12'sd-1370, 13'sd2551}},
{{12'sd2013, 13'sd2630, 12'sd-1835}, {12'sd-1886, 12'sd-2020, 11'sd-825}, {11'sd-887, 12'sd1329, 12'sd1999}},
{{12'sd1883, 13'sd2306, 12'sd-1270}, {11'sd-651, 13'sd-2266, 13'sd-2048}, {11'sd609, 11'sd-678, 13'sd-2530}},
{{13'sd2068, 11'sd991, 10'sd-258}, {12'sd-1826, 10'sd-496, 13'sd2668}, {12'sd1374, 12'sd-1934, 13'sd3269}},
{{8'sd66, 11'sd948, 11'sd-519}, {13'sd2270, 13'sd-2771, 9'sd245}, {12'sd1397, 13'sd-2233, 9'sd231}},
{{10'sd379, 12'sd-1518, 10'sd-489}, {11'sd-989, 12'sd1884, 12'sd-1593}, {11'sd-525, 12'sd-1870, 10'sd258}},
{{11'sd990, 12'sd1696, 12'sd1716}, {12'sd1593, 12'sd-1835, 12'sd-1091}, {12'sd-1292, 13'sd-2243, 11'sd781}},
{{13'sd2116, 13'sd2639, 12'sd1875}, {12'sd-1259, 11'sd-736, 11'sd-875}, {13'sd2326, 11'sd861, 13'sd-2095}},
{{10'sd314, 10'sd-365, 12'sd-1568}, {10'sd-397, 12'sd1100, 13'sd-2148}, {13'sd-2286, 12'sd-2044, 13'sd2103}},
{{7'sd38, 10'sd362, 12'sd1391}, {12'sd1232, 12'sd-1744, 13'sd-2072}, {13'sd2600, 13'sd2291, 11'sd-739}},
{{11'sd575, 12'sd1492, 12'sd-1716}, {12'sd1079, 10'sd-315, 8'sd79}, {12'sd-1420, 12'sd1035, 12'sd-1671}},
{{13'sd2414, 12'sd1946, 11'sd557}, {11'sd-847, 12'sd-1993, 11'sd-800}, {13'sd2691, 12'sd-1035, 13'sd2297}},
{{9'sd172, 13'sd-2636, 13'sd-2304}, {12'sd1101, 12'sd1259, 10'sd471}, {13'sd-2419, 10'sd-342, 12'sd-1218}},
{{13'sd2489, 11'sd-668, 13'sd2428}, {12'sd1867, 13'sd-2410, 12'sd1514}, {12'sd1156, 12'sd1218, 14'sd-4275}},
{{11'sd997, 13'sd2071, 10'sd359}, {12'sd1899, 10'sd-506, 8'sd88}, {11'sd-886, 11'sd640, 10'sd302}},
{{11'sd660, 11'sd-964, 11'sd889}, {13'sd-2077, 11'sd885, 12'sd1311}, {12'sd1376, 10'sd352, 12'sd1719}},
{{12'sd-1267, 12'sd-1837, 12'sd-1774}, {13'sd-2426, 11'sd963, 13'sd2602}, {13'sd2068, 9'sd232, 12'sd1613}},
{{11'sd649, 13'sd-2171, 10'sd-498}, {12'sd1242, 3'sd-3, 12'sd1533}, {12'sd-1089, 13'sd2690, 12'sd-1268}},
{{12'sd-1595, 12'sd1175, 9'sd246}, {12'sd-1249, 13'sd3658, 12'sd1135}, {11'sd811, 12'sd-1677, 13'sd2820}},
{{11'sd932, 12'sd-1570, 13'sd2995}, {13'sd-2294, 9'sd-141, 12'sd1771}, {12'sd1408, 8'sd-102, 12'sd1757}},
{{12'sd1549, 9'sd-187, 8'sd-107}, {12'sd1575, 13'sd2456, 12'sd-1665}, {9'sd254, 12'sd1682, 13'sd2694}},
{{13'sd-2720, 12'sd-1361, 9'sd-215}, {12'sd-1784, 12'sd-1133, 11'sd656}, {12'sd1177, 7'sd54, 12'sd1475}},
{{12'sd-1226, 12'sd-1697, 11'sd-544}, {13'sd2564, 12'sd-1193, 11'sd824}, {13'sd2287, 9'sd129, 10'sd-490}},
{{8'sd75, 12'sd1345, 12'sd1450}, {13'sd2295, 12'sd1842, 8'sd-83}, {10'sd490, 13'sd2474, 10'sd-426}},
{{13'sd2851, 11'sd670, 11'sd-816}, {12'sd1136, 12'sd-1975, 12'sd-1727}, {12'sd-1608, 11'sd-979, 7'sd59}}},
{
{{12'sd1046, 10'sd-472, 13'sd2219}, {13'sd2402, 12'sd1627, 12'sd-1091}, {12'sd-1548, 12'sd-1672, 12'sd-1852}},
{{13'sd-2529, 13'sd-2225, 13'sd-3565}, {11'sd584, 10'sd-268, 10'sd-409}, {12'sd1299, 12'sd1617, 13'sd-3225}},
{{12'sd-1352, 6'sd27, 13'sd-4084}, {14'sd-4400, 12'sd-1108, 11'sd842}, {12'sd-1305, 13'sd3085, 10'sd-363}},
{{12'sd-1223, 13'sd2411, 13'sd-2366}, {11'sd-1005, 10'sd-275, 12'sd1198}, {9'sd-220, 11'sd896, 12'sd1073}},
{{12'sd-1202, 13'sd-2631, 8'sd-65}, {12'sd-1721, 10'sd-365, 11'sd528}, {10'sd480, 12'sd-1070, 12'sd1854}},
{{12'sd1867, 8'sd-89, 12'sd1349}, {12'sd1924, 11'sd687, 12'sd1157}, {12'sd1983, 12'sd1072, 12'sd1979}},
{{12'sd1211, 9'sd-189, 13'sd2353}, {12'sd1654, 13'sd-2333, 13'sd2767}, {12'sd-1571, 12'sd1464, 12'sd-1651}},
{{8'sd65, 13'sd2846, 10'sd405}, {13'sd2569, 12'sd-1647, 12'sd1554}, {9'sd242, 12'sd-1944, 12'sd-1957}},
{{11'sd694, 11'sd643, 12'sd-1881}, {13'sd-3415, 11'sd766, 12'sd-1175}, {11'sd760, 12'sd-1406, 13'sd-3941}},
{{13'sd-2784, 13'sd2453, 11'sd-579}, {13'sd-2702, 10'sd449, 11'sd-524}, {11'sd602, 11'sd600, 11'sd-600}},
{{13'sd3777, 10'sd390, 12'sd2007}, {12'sd1868, 8'sd-97, 12'sd-1181}, {11'sd-847, 12'sd-1631, 14'sd5029}},
{{10'sd-408, 11'sd663, 8'sd-79}, {12'sd-1205, 10'sd-374, 12'sd-1408}, {11'sd-615, 12'sd1621, 12'sd-1199}},
{{10'sd488, 12'sd-1744, 12'sd-1311}, {12'sd-1172, 12'sd1344, 12'sd-1233}, {13'sd3632, 13'sd3263, 12'sd1989}},
{{13'sd2921, 9'sd-203, 11'sd632}, {12'sd-1122, 12'sd-1864, 12'sd-1504}, {13'sd2428, 12'sd1494, 11'sd613}},
{{12'sd-1066, 12'sd-1168, 10'sd-279}, {11'sd640, 13'sd-2669, 12'sd-1799}, {13'sd2176, 12'sd1130, 11'sd682}},
{{12'sd1220, 12'sd-1428, 12'sd-1462}, {13'sd-2597, 13'sd2064, 7'sd-34}, {12'sd1765, 13'sd2397, 10'sd-492}},
{{13'sd2493, 12'sd1561, 10'sd502}, {10'sd466, 13'sd2283, 11'sd-904}, {13'sd2597, 12'sd-1581, 11'sd729}},
{{10'sd384, 11'sd-730, 7'sd-58}, {13'sd-2600, 11'sd-863, 13'sd-3124}, {12'sd1231, 13'sd2131, 12'sd-1122}},
{{12'sd-1098, 12'sd1830, 12'sd1344}, {13'sd2301, 9'sd-178, 11'sd715}, {10'sd262, 12'sd-2046, 12'sd-1817}},
{{11'sd602, 9'sd244, 11'sd963}, {11'sd-631, 8'sd-113, 12'sd-1292}, {11'sd-601, 12'sd1331, 12'sd1408}},
{{12'sd-1537, 11'sd-846, 13'sd-3414}, {13'sd-2742, 12'sd2006, 13'sd-2155}, {12'sd-1344, 13'sd-2268, 12'sd-1116}},
{{13'sd-2434, 11'sd-934, 11'sd-738}, {12'sd-1683, 12'sd1293, 11'sd-650}, {11'sd767, 11'sd-840, 12'sd-1827}},
{{8'sd106, 10'sd-347, 12'sd1932}, {11'sd512, 13'sd-2433, 12'sd1824}, {10'sd-510, 11'sd-883, 12'sd-1295}},
{{8'sd-104, 12'sd1168, 11'sd-565}, {13'sd-2908, 13'sd2160, 12'sd1301}, {12'sd-1890, 12'sd-2029, 12'sd1810}},
{{13'sd-3584, 11'sd640, 12'sd-1275}, {13'sd-2532, 9'sd-235, 13'sd-2464}, {12'sd-1029, 13'sd-3581, 12'sd-2021}},
{{12'sd1610, 12'sd-1987, 13'sd-2834}, {9'sd-169, 12'sd1178, 12'sd1292}, {11'sd-756, 10'sd-308, 13'sd2251}},
{{10'sd-280, 10'sd357, 13'sd-2091}, {11'sd-687, 12'sd-1954, 12'sd-1301}, {13'sd-2726, 9'sd-205, 9'sd236}},
{{8'sd-91, 7'sd-43, 10'sd501}, {12'sd-1884, 13'sd-2135, 12'sd1793}, {9'sd-199, 13'sd2191, 12'sd-1541}},
{{11'sd966, 13'sd-2818, 13'sd-3134}, {12'sd-1120, 12'sd1474, 11'sd885}, {12'sd-1884, 12'sd1478, 8'sd115}},
{{13'sd-3797, 9'sd-199, 12'sd-1105}, {10'sd-373, 13'sd2096, 10'sd-278}, {13'sd2614, 13'sd2416, 13'sd3068}},
{{11'sd-910, 12'sd-1397, 9'sd-213}, {12'sd-1511, 11'sd780, 12'sd-1758}, {12'sd1290, 13'sd-2658, 10'sd-409}},
{{13'sd3950, 13'sd3514, 12'sd-1747}, {10'sd-278, 13'sd3510, 12'sd1358}, {10'sd-404, 11'sd900, 12'sd-1913}},
{{8'sd-113, 13'sd-2323, 11'sd-891}, {12'sd1710, 13'sd2616, 12'sd1786}, {13'sd-2329, 11'sd740, 12'sd-1434}},
{{13'sd-3077, 12'sd-1689, 7'sd-40}, {12'sd-1968, 8'sd-81, 12'sd-1364}, {13'sd2626, 11'sd-800, 12'sd-1299}},
{{13'sd2282, 12'sd2028, 13'sd2641}, {12'sd-1279, 10'sd324, 11'sd-643}, {13'sd2438, 13'sd-2129, 11'sd593}},
{{12'sd-1200, 12'sd-1324, 11'sd-590}, {11'sd541, 11'sd-763, 11'sd916}, {12'sd-1906, 12'sd-1387, 10'sd-511}},
{{12'sd1797, 12'sd1526, 11'sd-533}, {13'sd-2830, 12'sd1128, 13'sd-2284}, {11'sd-997, 12'sd1739, 13'sd2087}},
{{12'sd1342, 13'sd2157, 12'sd1595}, {12'sd1269, 13'sd2688, 9'sd-169}, {12'sd1934, 11'sd519, 13'sd-2048}},
{{12'sd1240, 11'sd-537, 13'sd-3089}, {9'sd252, 13'sd-2069, 11'sd535}, {12'sd1339, 12'sd1251, 10'sd446}},
{{10'sd-381, 12'sd1906, 13'sd2747}, {13'sd-2196, 12'sd-1722, 13'sd-2161}, {5'sd-8, 12'sd-1606, 11'sd-816}},
{{12'sd-1079, 13'sd2334, 11'sd-869}, {13'sd2496, 13'sd-2193, 12'sd1730}, {11'sd-596, 12'sd1988, 12'sd1751}},
{{12'sd1228, 13'sd2925, 12'sd-1489}, {12'sd-1658, 12'sd1605, 12'sd-1679}, {13'sd-3002, 10'sd305, 13'sd-2397}},
{{12'sd1457, 12'sd-1701, 10'sd312}, {12'sd1178, 7'sd-43, 7'sd-32}, {10'sd430, 9'sd213, 11'sd815}},
{{12'sd1990, 13'sd-2297, 13'sd2242}, {13'sd-2277, 13'sd-2775, 6'sd-26}, {13'sd2961, 9'sd208, 13'sd2936}},
{{10'sd-346, 9'sd153, 10'sd-409}, {13'sd-2182, 7'sd47, 13'sd-2076}, {13'sd2155, 13'sd-2486, 10'sd-306}},
{{12'sd-1828, 12'sd-1658, 11'sd991}, {9'sd252, 11'sd686, 11'sd-912}, {13'sd-3272, 12'sd-1712, 12'sd-1260}},
{{9'sd-191, 12'sd1390, 13'sd-2396}, {10'sd479, 13'sd2495, 10'sd-439}, {11'sd-530, 13'sd2307, 12'sd-1570}},
{{10'sd-391, 13'sd-2404, 12'sd1079}, {12'sd-1771, 12'sd-1748, 12'sd-1362}, {13'sd-2769, 10'sd277, 10'sd320}},
{{12'sd1186, 11'sd-606, 7'sd42}, {10'sd347, 13'sd-2198, 7'sd-53}, {13'sd2613, 7'sd-50, 12'sd-1990}},
{{10'sd323, 13'sd-2184, 12'sd1777}, {13'sd2342, 11'sd-914, 10'sd498}, {12'sd1428, 7'sd51, 12'sd1481}},
{{12'sd-1258, 13'sd-2461, 12'sd-1092}, {12'sd1233, 12'sd-1566, 11'sd-838}, {12'sd-1785, 12'sd1087, 12'sd-1345}},
{{13'sd-2217, 13'sd-2281, 12'sd1999}, {13'sd-2217, 11'sd665, 8'sd113}, {13'sd2823, 10'sd-366, 12'sd-1141}},
{{12'sd-1862, 13'sd2195, 14'sd4700}, {5'sd-13, 12'sd-1545, 12'sd1578}, {13'sd-3918, 11'sd-688, 11'sd-550}},
{{12'sd1073, 12'sd1030, 12'sd-1431}, {12'sd-1350, 11'sd619, 10'sd-316}, {12'sd-1276, 13'sd2201, 11'sd-628}},
{{12'sd1819, 12'sd-1266, 12'sd-1531}, {13'sd-2515, 11'sd724, 12'sd1754}, {11'sd-779, 12'sd1307, 10'sd-402}},
{{11'sd-556, 5'sd14, 12'sd-1625}, {11'sd-788, 12'sd1425, 12'sd1137}, {13'sd2279, 13'sd2571, 10'sd340}},
{{13'sd-2842, 12'sd1179, 12'sd-1255}, {13'sd-3021, 12'sd2033, 13'sd-3036}, {12'sd1971, 12'sd1188, 10'sd-412}},
{{14'sd4375, 12'sd1536, 12'sd-1674}, {13'sd2981, 8'sd124, 10'sd-434}, {12'sd-1479, 13'sd2912, 13'sd-2990}},
{{13'sd4062, 11'sd646, 13'sd-3195}, {14'sd5021, 12'sd-1777, 12'sd1244}, {9'sd163, 13'sd2445, 9'sd-163}},
{{11'sd-662, 12'sd-1202, 11'sd-798}, {11'sd949, 10'sd383, 12'sd1704}, {11'sd-701, 10'sd469, 11'sd-952}},
{{11'sd922, 13'sd2644, 12'sd-1505}, {13'sd2321, 13'sd3329, 10'sd261}, {6'sd20, 11'sd881, 13'sd-2466}},
{{12'sd1702, 12'sd1966, 12'sd1910}, {12'sd1071, 12'sd1381, 12'sd1695}, {12'sd1826, 12'sd-2005, 12'sd-1662}},
{{11'sd802, 13'sd-2305, 11'sd812}, {13'sd2586, 12'sd1509, 12'sd-1714}, {10'sd480, 13'sd-2400, 12'sd-1409}},
{{12'sd1066, 12'sd-1571, 10'sd316}, {10'sd-269, 12'sd-1370, 10'sd264}, {12'sd-1227, 12'sd1269, 13'sd-2292}}},
{
{{12'sd1223, 12'sd-1069, 7'sd53}, {13'sd2196, 13'sd3199, 8'sd-90}, {11'sd-793, 13'sd2528, 13'sd-2168}},
{{9'sd195, 11'sd672, 12'sd1532}, {12'sd1548, 12'sd1299, 11'sd613}, {10'sd-459, 13'sd2445, 9'sd-248}},
{{13'sd-2280, 13'sd-2518, 13'sd-2457}, {13'sd2587, 9'sd187, 8'sd110}, {13'sd2315, 8'sd-84, 13'sd2338}},
{{13'sd-2854, 12'sd-1996, 12'sd1334}, {12'sd-1510, 11'sd-646, 11'sd-717}, {11'sd787, 13'sd2788, 12'sd-1099}},
{{13'sd-2053, 11'sd-526, 13'sd-2684}, {13'sd-2166, 12'sd1164, 12'sd1528}, {10'sd314, 12'sd1409, 12'sd-2024}},
{{11'sd584, 13'sd2540, 11'sd-1003}, {13'sd2324, 13'sd2069, 12'sd1157}, {11'sd-543, 13'sd2143, 11'sd-760}},
{{13'sd2074, 10'sd-317, 12'sd-1731}, {13'sd-3036, 13'sd-2315, 12'sd1910}, {13'sd-2310, 12'sd-1323, 12'sd-1396}},
{{12'sd-1975, 11'sd745, 12'sd-1942}, {13'sd2608, 12'sd-1408, 13'sd2559}, {11'sd908, 11'sd667, 12'sd1783}},
{{11'sd-780, 12'sd-1849, 11'sd775}, {12'sd1378, 12'sd-1210, 13'sd-2058}, {13'sd-2189, 8'sd-81, 13'sd2130}},
{{9'sd181, 11'sd1002, 11'sd-718}, {12'sd1984, 9'sd-215, 13'sd-2760}, {12'sd-1937, 13'sd2610, 11'sd777}},
{{13'sd2651, 9'sd-177, 14'sd4760}, {12'sd-1676, 13'sd2857, 12'sd-1328}, {12'sd1530, 13'sd3368, 11'sd-657}},
{{12'sd1365, 10'sd500, 12'sd1696}, {12'sd-1571, 11'sd-783, 13'sd2791}, {13'sd2221, 12'sd1129, 12'sd-1182}},
{{13'sd-2445, 12'sd-2026, 14'sd-4705}, {12'sd1955, 13'sd-2340, 13'sd-3223}, {12'sd-1370, 12'sd-1117, 11'sd-573}},
{{12'sd-1059, 12'sd-1936, 10'sd485}, {13'sd-2454, 11'sd-782, 12'sd1715}, {12'sd1437, 11'sd777, 13'sd2620}},
{{12'sd1765, 10'sd-476, 12'sd-1735}, {10'sd-415, 13'sd2400, 13'sd2224}, {12'sd-1430, 12'sd1437, 13'sd-2715}},
{{11'sd-846, 13'sd2162, 12'sd-1158}, {13'sd-2101, 12'sd-1671, 13'sd-2566}, {11'sd-534, 7'sd32, 10'sd-424}},
{{13'sd-2057, 11'sd-539, 13'sd-2836}, {9'sd-129, 13'sd2754, 11'sd-656}, {10'sd-372, 13'sd-2370, 12'sd-1684}},
{{12'sd1260, 12'sd1258, 13'sd-2575}, {12'sd1224, 12'sd1258, 13'sd-2234}, {13'sd2991, 12'sd1765, 12'sd1190}},
{{12'sd1321, 13'sd2583, 11'sd890}, {9'sd-216, 12'sd1073, 13'sd2345}, {10'sd-435, 13'sd2473, 11'sd-541}},
{{13'sd-2065, 12'sd-1222, 9'sd-224}, {12'sd-1967, 11'sd917, 13'sd-3211}, {9'sd132, 10'sd324, 9'sd195}},
{{12'sd1467, 10'sd-263, 12'sd1392}, {13'sd-2684, 13'sd-2447, 12'sd-1819}, {10'sd-334, 10'sd-436, 12'sd-1726}},
{{13'sd-3073, 8'sd-119, 13'sd3545}, {11'sd-609, 13'sd-3666, 9'sd153}, {11'sd732, 12'sd1589, 12'sd1567}},
{{13'sd-2558, 11'sd-802, 13'sd2232}, {13'sd2847, 13'sd2484, 12'sd-1304}, {11'sd-920, 11'sd-895, 13'sd-2906}},
{{10'sd386, 12'sd1826, 13'sd-2597}, {12'sd-1857, 13'sd-2855, 12'sd1717}, {12'sd1678, 13'sd2179, 12'sd-1583}},
{{8'sd81, 13'sd-2418, 10'sd408}, {13'sd2500, 10'sd351, 9'sd-247}, {13'sd-2159, 13'sd-3128, 11'sd526}},
{{10'sd-484, 12'sd1577, 12'sd-1149}, {12'sd-1244, 11'sd-684, 13'sd2504}, {11'sd997, 10'sd-264, 12'sd1416}},
{{12'sd1666, 13'sd-2312, 12'sd-1203}, {11'sd-676, 13'sd-2253, 13'sd2880}, {8'sd-84, 12'sd1053, 12'sd1884}},
{{12'sd1597, 12'sd1152, 12'sd1426}, {13'sd2327, 11'sd-636, 12'sd-1621}, {10'sd507, 12'sd1771, 13'sd2532}},
{{13'sd-2918, 11'sd535, 12'sd2027}, {12'sd1081, 4'sd-7, 13'sd-2080}, {10'sd366, 12'sd-1225, 12'sd1654}},
{{12'sd-1427, 10'sd-323, 13'sd3567}, {13'sd-3929, 13'sd-2775, 12'sd-1298}, {11'sd795, 12'sd1155, 11'sd-828}},
{{13'sd2295, 13'sd-2065, 12'sd1960}, {12'sd1742, 5'sd-10, 12'sd1862}, {13'sd2431, 12'sd1382, 13'sd-2251}},
{{12'sd-1580, 13'sd3725, 8'sd-119}, {12'sd1100, 10'sd-363, 12'sd-1563}, {11'sd-904, 13'sd2555, 13'sd2614}},
{{11'sd-912, 11'sd-972, 12'sd1907}, {13'sd2906, 10'sd-497, 12'sd-1546}, {13'sd2454, 12'sd-1904, 10'sd266}},
{{11'sd-796, 11'sd869, 13'sd2366}, {12'sd-1517, 12'sd-1748, 12'sd-1969}, {12'sd-1989, 12'sd1135, 11'sd512}},
{{11'sd784, 12'sd1268, 10'sd-401}, {11'sd844, 12'sd1178, 11'sd849}, {12'sd-1410, 13'sd2054, 12'sd1985}},
{{12'sd-1939, 13'sd-2474, 12'sd-1451}, {13'sd2387, 12'sd1480, 9'sd205}, {12'sd-1699, 12'sd1989, 12'sd-1952}},
{{13'sd-2478, 12'sd-1803, 11'sd651}, {12'sd-1337, 12'sd1883, 11'sd-586}, {12'sd1072, 12'sd1964, 12'sd1323}},
{{12'sd-1848, 9'sd-142, 10'sd-322}, {12'sd-1364, 13'sd3386, 12'sd1110}, {13'sd-2840, 13'sd-2086, 10'sd475}},
{{12'sd-1929, 12'sd-1457, 14'sd-4537}, {9'sd133, 11'sd929, 11'sd-520}, {13'sd2376, 11'sd617, 13'sd-2599}},
{{9'sd-173, 11'sd518, 13'sd-2329}, {12'sd1144, 12'sd1458, 12'sd2018}, {13'sd2821, 12'sd-1778, 11'sd603}},
{{11'sd649, 13'sd-2501, 10'sd358}, {3'sd3, 10'sd-484, 12'sd-1040}, {11'sd764, 13'sd-3358, 11'sd-513}},
{{10'sd-471, 12'sd1076, 12'sd-1536}, {13'sd-2901, 12'sd1600, 12'sd1368}, {12'sd-1106, 10'sd-266, 12'sd-1194}},
{{12'sd1532, 13'sd2471, 13'sd2381}, {10'sd481, 11'sd572, 12'sd1837}, {13'sd-2373, 6'sd16, 13'sd-2720}},
{{13'sd2847, 10'sd413, 12'sd1243}, {10'sd443, 13'sd-2674, 11'sd965}, {13'sd-2986, 10'sd482, 12'sd-1729}},
{{11'sd831, 12'sd-1578, 12'sd1840}, {9'sd-200, 11'sd-646, 6'sd18}, {13'sd2153, 11'sd869, 12'sd-1293}},
{{12'sd-1882, 12'sd-1504, 13'sd-3441}, {4'sd4, 9'sd-222, 12'sd-1453}, {12'sd1906, 10'sd-469, 12'sd-2025}},
{{13'sd2143, 12'sd1470, 12'sd1427}, {13'sd2432, 11'sd741, 12'sd-1068}, {11'sd562, 13'sd2462, 12'sd1866}},
{{13'sd2128, 12'sd-2019, 13'sd-2087}, {11'sd994, 12'sd-1024, 12'sd-1909}, {6'sd-29, 12'sd-1675, 11'sd993}},
{{12'sd-1516, 12'sd1349, 9'sd-239}, {11'sd681, 11'sd-881, 13'sd2075}, {13'sd-2433, 10'sd-415, 13'sd2478}},
{{11'sd-743, 12'sd1492, 11'sd792}, {13'sd-2860, 13'sd-2234, 11'sd825}, {13'sd-2681, 12'sd1060, 11'sd550}},
{{12'sd-1669, 11'sd-517, 12'sd1168}, {13'sd-2744, 13'sd2244, 13'sd2827}, {11'sd-561, 12'sd-1363, 10'sd433}},
{{13'sd2305, 12'sd-1495, 11'sd-612}, {13'sd-2411, 12'sd1201, 12'sd1734}, {11'sd654, 11'sd891, 13'sd2993}},
{{13'sd-2221, 12'sd-1133, 9'sd176}, {13'sd-3479, 13'sd-2146, 11'sd855}, {12'sd-1656, 12'sd1258, 13'sd2453}},
{{9'sd237, 12'sd1503, 13'sd-3023}, {12'sd1911, 13'sd2740, 13'sd-2882}, {12'sd1858, 11'sd-572, 13'sd-2054}},
{{13'sd2331, 11'sd767, 11'sd742}, {12'sd1707, 10'sd256, 10'sd471}, {11'sd-939, 13'sd-2693, 12'sd1330}},
{{13'sd2679, 13'sd2651, 8'sd94}, {13'sd2737, 12'sd-1710, 11'sd-881}, {12'sd1196, 8'sd-81, 11'sd-983}},
{{13'sd-2627, 12'sd1525, 13'sd-2440}, {10'sd424, 12'sd1425, 12'sd2005}, {6'sd-18, 11'sd569, 13'sd-3018}},
{{13'sd3799, 11'sd-602, 13'sd-3553}, {13'sd2130, 12'sd1101, 12'sd-1373}, {13'sd3090, 13'sd3365, 13'sd2773}},
{{13'sd2923, 11'sd611, 12'sd1345}, {12'sd2043, 11'sd-786, 12'sd-1619}, {14'sd4732, 9'sd215, 10'sd-319}},
{{12'sd-1473, 10'sd392, 12'sd-1796}, {13'sd-2781, 10'sd-416, 11'sd-793}, {12'sd1978, 13'sd2766, 11'sd-577}},
{{11'sd-537, 13'sd-2491, 12'sd-1268}, {12'sd1960, 9'sd-241, 13'sd-2081}, {12'sd-1101, 13'sd2140, 13'sd-3153}},
{{11'sd-929, 12'sd1053, 10'sd-349}, {12'sd1803, 9'sd-226, 13'sd2625}, {10'sd417, 12'sd1812, 12'sd-2001}},
{{12'sd1589, 11'sd-771, 10'sd316}, {13'sd-2415, 12'sd-1548, 12'sd1413}, {12'sd-1469, 11'sd-541, 11'sd-1014}},
{{12'sd-1160, 12'sd-1207, 11'sd-677}, {12'sd-1239, 13'sd2129, 11'sd-815}, {13'sd-2427, 12'sd-1631, 12'sd1915}}},
{
{{12'sd-1881, 12'sd-1304, 12'sd-1435}, {13'sd3196, 12'sd-1884, 13'sd3005}, {9'sd-145, 10'sd426, 12'sd-1599}},
{{12'sd-1836, 11'sd-743, 12'sd1908}, {13'sd-2095, 11'sd-627, 11'sd-622}, {9'sd-194, 11'sd561, 13'sd-2570}},
{{13'sd3159, 13'sd3455, 9'sd233}, {13'sd2693, 13'sd2684, 11'sd-513}, {13'sd2380, 8'sd-99, 13'sd-2777}},
{{13'sd-2339, 13'sd-2758, 12'sd1050}, {12'sd-1362, 11'sd-722, 12'sd-1244}, {12'sd-1623, 13'sd-2661, 12'sd1719}},
{{12'sd-1221, 12'sd-1885, 12'sd1948}, {12'sd1514, 13'sd-2602, 11'sd714}, {10'sd280, 10'sd-303, 9'sd-155}},
{{9'sd238, 11'sd849, 12'sd2019}, {9'sd218, 12'sd1193, 10'sd318}, {9'sd-231, 10'sd330, 12'sd2021}},
{{13'sd-2735, 11'sd681, 10'sd411}, {13'sd2080, 13'sd-2161, 12'sd-2029}, {13'sd2443, 13'sd-2271, 12'sd-2043}},
{{13'sd-2991, 11'sd-542, 12'sd-1170}, {13'sd-2134, 11'sd758, 11'sd601}, {13'sd2630, 13'sd-2290, 10'sd-313}},
{{12'sd1941, 12'sd1643, 8'sd96}, {12'sd-2016, 11'sd-778, 12'sd1353}, {13'sd-2096, 13'sd2233, 12'sd1657}},
{{13'sd2679, 13'sd2712, 9'sd151}, {8'sd101, 10'sd-298, 13'sd2277}, {11'sd656, 13'sd-2399, 12'sd-1099}},
{{12'sd-1880, 9'sd156, 13'sd2363}, {13'sd-3457, 13'sd-2630, 8'sd74}, {13'sd-2984, 13'sd-2696, 12'sd-1851}},
{{11'sd678, 12'sd-1944, 13'sd2352}, {10'sd303, 11'sd-597, 12'sd1389}, {9'sd191, 12'sd-1133, 9'sd-140}},
{{13'sd-2642, 13'sd2238, 10'sd389}, {12'sd-1144, 11'sd590, 12'sd1350}, {13'sd3073, 12'sd-1761, 13'sd-2469}},
{{13'sd-2426, 11'sd931, 13'sd2429}, {10'sd308, 13'sd-2839, 12'sd1899}, {12'sd-1457, 11'sd-578, 12'sd1929}},
{{13'sd-2302, 11'sd-575, 11'sd552}, {9'sd-199, 10'sd-277, 11'sd662}, {12'sd1734, 12'sd1304, 10'sd483}},
{{10'sd269, 12'sd-1228, 12'sd1467}, {12'sd-1423, 12'sd-1190, 12'sd1238}, {10'sd-386, 12'sd1444, 12'sd1919}},
{{13'sd2181, 13'sd-2980, 13'sd-3211}, {13'sd2617, 8'sd112, 12'sd-1325}, {12'sd1566, 10'sd371, 11'sd514}},
{{7'sd-60, 12'sd-1458, 13'sd2800}, {12'sd-1985, 12'sd1740, 12'sd1548}, {13'sd-2830, 10'sd443, 11'sd-936}},
{{12'sd1906, 12'sd-1344, 11'sd-1020}, {13'sd2910, 10'sd471, 12'sd1879}, {13'sd2157, 12'sd1205, 9'sd189}},
{{12'sd-1956, 10'sd-479, 11'sd915}, {10'sd-430, 12'sd2046, 12'sd1907}, {12'sd-1265, 12'sd-1403, 11'sd-995}},
{{13'sd2373, 9'sd-184, 12'sd1349}, {13'sd-2447, 13'sd-2346, 12'sd1479}, {13'sd-3189, 11'sd-821, 12'sd-1137}},
{{11'sd1002, 13'sd-2697, 13'sd2294}, {6'sd31, 13'sd-2393, 13'sd-2405}, {13'sd-2659, 13'sd-2068, 11'sd572}},
{{13'sd2767, 10'sd436, 12'sd1856}, {13'sd-2129, 12'sd-1175, 10'sd256}, {9'sd221, 12'sd-1295, 12'sd-1937}},
{{12'sd-1834, 12'sd-1092, 10'sd299}, {12'sd1399, 12'sd-1237, 12'sd-1478}, {13'sd-2144, 10'sd-346, 9'sd-195}},
{{14'sd4214, 14'sd4585, 13'sd2469}, {7'sd-40, 12'sd1617, 9'sd-195}, {12'sd1624, 7'sd-42, 10'sd-398}},
{{12'sd1479, 13'sd-2561, 13'sd-2419}, {13'sd2603, 13'sd2558, 12'sd-1920}, {11'sd880, 13'sd2663, 10'sd-489}},
{{12'sd-1516, 12'sd1920, 12'sd-1457}, {8'sd-125, 10'sd-294, 10'sd286}, {6'sd-26, 13'sd-2283, 12'sd-1899}},
{{11'sd842, 13'sd2623, 13'sd2415}, {8'sd-88, 13'sd2388, 13'sd2858}, {11'sd-934, 9'sd173, 12'sd-1647}},
{{13'sd-2339, 12'sd-1691, 12'sd-2013}, {13'sd-2827, 13'sd-2268, 12'sd-1413}, {12'sd1599, 12'sd1941, 11'sd-762}},
{{13'sd-2565, 12'sd-1789, 11'sd530}, {13'sd-2686, 9'sd138, 12'sd-1919}, {12'sd1355, 9'sd-179, 9'sd-219}},
{{12'sd1227, 12'sd1725, 12'sd-1728}, {13'sd-2349, 10'sd-286, 12'sd-1324}, {13'sd-2324, 11'sd554, 10'sd-387}},
{{10'sd-410, 12'sd-1311, 7'sd-47}, {12'sd1154, 13'sd2621, 11'sd857}, {9'sd-167, 11'sd-962, 12'sd1270}},
{{11'sd820, 13'sd-2385, 9'sd234}, {13'sd-2543, 10'sd-432, 12'sd-1686}, {10'sd-266, 12'sd1705, 13'sd-2940}},
{{12'sd1571, 8'sd-86, 12'sd-1145}, {12'sd1839, 13'sd-2083, 12'sd-1268}, {13'sd-2496, 12'sd1944, 13'sd-2340}},
{{9'sd-129, 12'sd-1806, 13'sd-2269}, {10'sd417, 12'sd-1432, 12'sd-1402}, {12'sd-1898, 12'sd-1040, 12'sd-1744}},
{{12'sd-1872, 12'sd1130, 12'sd1795}, {12'sd1296, 12'sd-1771, 10'sd-487}, {12'sd1994, 11'sd-890, 11'sd-605}},
{{12'sd-1838, 13'sd2085, 13'sd2668}, {12'sd-1381, 6'sd17, 10'sd284}, {10'sd401, 12'sd1722, 10'sd-445}},
{{11'sd-711, 11'sd-585, 11'sd749}, {9'sd209, 13'sd-2541, 13'sd3622}, {10'sd330, 11'sd-747, 12'sd1564}},
{{12'sd-1836, 13'sd-2307, 13'sd-3073}, {12'sd1455, 13'sd-2048, 13'sd-2284}, {4'sd4, 10'sd484, 9'sd145}},
{{12'sd-1072, 11'sd-756, 12'sd1485}, {13'sd2457, 13'sd2268, 13'sd2106}, {10'sd-288, 12'sd1556, 10'sd-494}},
{{8'sd-107, 13'sd2971, 13'sd-3264}, {11'sd1009, 11'sd860, 10'sd333}, {12'sd-1868, 13'sd-2143, 12'sd-1675}},
{{13'sd2717, 13'sd2078, 13'sd2272}, {12'sd2017, 12'sd1663, 9'sd132}, {13'sd3035, 12'sd-1566, 11'sd896}},
{{12'sd-1091, 13'sd-2139, 12'sd1488}, {13'sd-2120, 9'sd171, 11'sd821}, {12'sd1356, 12'sd1370, 11'sd-828}},
{{11'sd835, 13'sd2308, 13'sd-2412}, {12'sd-1649, 10'sd502, 12'sd-1629}, {10'sd-435, 12'sd1944, 8'sd69}},
{{12'sd-1186, 12'sd1847, 12'sd-1190}, {12'sd1292, 13'sd-2703, 12'sd1610}, {12'sd-2026, 12'sd-1553, 10'sd356}},
{{12'sd2031, 12'sd1504, 11'sd925}, {13'sd-3129, 13'sd-2131, 11'sd763}, {11'sd-794, 11'sd897, 13'sd-2713}},
{{11'sd1006, 12'sd1834, 11'sd-601}, {11'sd995, 13'sd-2507, 11'sd-520}, {11'sd-634, 12'sd-1579, 12'sd1806}},
{{12'sd-1930, 9'sd230, 12'sd1795}, {11'sd-666, 12'sd-1419, 12'sd-2016}, {13'sd-2299, 10'sd293, 10'sd-477}},
{{13'sd-2073, 13'sd-2625, 12'sd-1829}, {11'sd-726, 13'sd2630, 10'sd304}, {13'sd2513, 11'sd572, 12'sd1031}},
{{8'sd80, 12'sd-1773, 9'sd252}, {13'sd2156, 12'sd1876, 13'sd2534}, {13'sd2128, 11'sd-963, 13'sd2973}},
{{4'sd-7, 11'sd667, 10'sd-370}, {12'sd-1714, 11'sd-700, 12'sd1193}, {11'sd1002, 8'sd105, 12'sd1849}},
{{12'sd1946, 12'sd-1237, 12'sd1296}, {12'sd1540, 12'sd-1947, 12'sd-1529}, {12'sd1449, 10'sd318, 12'sd-1815}},
{{12'sd1781, 9'sd212, 12'sd-1092}, {12'sd-1677, 12'sd1291, 11'sd-670}, {11'sd740, 12'sd-1353, 13'sd2841}},
{{13'sd2743, 13'sd2320, 13'sd2413}, {12'sd-1761, 13'sd2341, 10'sd-264}, {9'sd-236, 12'sd1337, 13'sd-2922}},
{{11'sd626, 13'sd-2479, 13'sd2177}, {12'sd1357, 8'sd68, 12'sd-1232}, {13'sd2072, 11'sd-677, 11'sd-705}},
{{12'sd1680, 12'sd-1124, 13'sd2825}, {13'sd-2432, 12'sd-1088, 12'sd-1184}, {10'sd-267, 12'sd1945, 12'sd-2047}},
{{11'sd813, 11'sd672, 11'sd-666}, {13'sd-2798, 12'sd-1337, 11'sd808}, {12'sd1550, 13'sd-2349, 12'sd-1557}},
{{12'sd1678, 10'sd393, 11'sd-998}, {11'sd686, 12'sd1289, 12'sd-1641}, {11'sd928, 12'sd1082, 12'sd1993}},
{{12'sd-1691, 12'sd-1116, 13'sd2484}, {9'sd239, 11'sd-676, 12'sd-1815}, {12'sd-1751, 11'sd606, 10'sd339}},
{{13'sd-2672, 11'sd909, 11'sd-638}, {13'sd2550, 12'sd1574, 8'sd101}, {12'sd1765, 11'sd547, 10'sd-309}},
{{12'sd1283, 12'sd1553, 12'sd-1510}, {13'sd3181, 12'sd-1107, 11'sd-523}, {13'sd2131, 13'sd-2429, 13'sd2076}},
{{12'sd1147, 13'sd-2389, 12'sd1620}, {12'sd-1367, 13'sd2220, 12'sd-1343}, {10'sd494, 12'sd-1254, 11'sd919}},
{{13'sd2518, 13'sd2070, 11'sd-882}, {12'sd1772, 13'sd2737, 12'sd-1495}, {12'sd-1939, 13'sd2566, 11'sd-693}},
{{10'sd-266, 11'sd-835, 12'sd-1393}, {7'sd-33, 10'sd-429, 13'sd2955}, {13'sd2750, 10'sd-425, 13'sd3138}}}},
// Weights for conv4_weight
{
{
{{11'sd-521, 11'sd944, 13'sd-2592}, {13'sd-2855, 12'sd2020, 11'sd-793}, {11'sd-607, 11'sd563, 12'sd1552}},
{{12'sd2013, 11'sd663, 10'sd263}, {13'sd2592, 12'sd-1512, 13'sd-2578}, {12'sd-1477, 10'sd-452, 13'sd2593}},
{{11'sd-984, 8'sd111, 12'sd-1904}, {11'sd-653, 12'sd-1965, 12'sd-1724}, {13'sd2192, 13'sd2963, 12'sd-1036}},
{{9'sd-134, 13'sd2736, 12'sd1225}, {12'sd-1067, 11'sd961, 13'sd2050}, {12'sd1283, 11'sd900, 13'sd-2798}},
{{11'sd527, 10'sd480, 13'sd-2662}, {12'sd1201, 12'sd1763, 12'sd-1344}, {13'sd-2671, 9'sd201, 10'sd336}},
{{11'sd875, 11'sd-812, 10'sd367}, {11'sd543, 11'sd-756, 11'sd533}, {12'sd1088, 13'sd2447, 11'sd538}},
{{12'sd1740, 11'sd-859, 12'sd1473}, {11'sd-679, 9'sd-188, 12'sd1263}, {13'sd-3398, 7'sd-38, 12'sd1756}},
{{10'sd409, 11'sd-858, 13'sd2543}, {11'sd520, 10'sd452, 12'sd1248}, {13'sd-3058, 12'sd-1620, 10'sd-344}},
{{11'sd569, 10'sd326, 11'sd-723}, {11'sd-842, 12'sd-1985, 12'sd-1634}, {12'sd-1814, 13'sd-2148, 11'sd968}},
{{8'sd-87, 13'sd2060, 12'sd-1385}, {12'sd-1579, 13'sd2276, 13'sd-2160}, {11'sd896, 9'sd-151, 12'sd-1564}},
{{10'sd-455, 5'sd-14, 13'sd2418}, {9'sd-232, 12'sd1723, 12'sd-1717}, {12'sd-1495, 13'sd2943, 13'sd2296}},
{{12'sd-1865, 13'sd-2203, 12'sd-1935}, {5'sd-14, 11'sd-969, 13'sd2560}, {9'sd-129, 13'sd-2724, 13'sd-2361}},
{{12'sd1919, 11'sd-996, 11'sd-846}, {9'sd-151, 9'sd-160, 9'sd235}, {10'sd-327, 13'sd-2575, 12'sd-1424}},
{{12'sd-1397, 13'sd2377, 12'sd-1614}, {12'sd1061, 12'sd1554, 13'sd2220}, {10'sd349, 11'sd965, 13'sd-2479}},
{{11'sd513, 11'sd-962, 12'sd-1916}, {12'sd1086, 10'sd-366, 10'sd498}, {9'sd206, 10'sd-273, 12'sd-1320}},
{{7'sd-47, 12'sd1579, 9'sd143}, {13'sd2502, 11'sd-1022, 12'sd-1884}, {11'sd-616, 12'sd1471, 13'sd-2240}},
{{13'sd-3146, 12'sd-1369, 12'sd-1327}, {12'sd1571, 12'sd-1379, 13'sd-2627}, {11'sd-851, 11'sd605, 13'sd-2915}},
{{11'sd-604, 13'sd2746, 10'sd405}, {13'sd2325, 13'sd3207, 11'sd-558}, {12'sd-1624, 13'sd2095, 12'sd1540}},
{{13'sd2939, 11'sd-764, 12'sd1771}, {13'sd-2416, 13'sd-2884, 12'sd1922}, {12'sd1455, 11'sd-524, 12'sd2019}},
{{11'sd826, 13'sd3047, 13'sd3006}, {10'sd-441, 12'sd1861, 12'sd-1327}, {11'sd876, 12'sd-1073, 10'sd-313}},
{{12'sd-1239, 12'sd-1041, 10'sd-269}, {11'sd-782, 13'sd-2317, 13'sd-2557}, {12'sd1355, 13'sd-2244, 13'sd-3073}},
{{13'sd-2140, 9'sd233, 10'sd-424}, {13'sd-2445, 12'sd1286, 12'sd1923}, {12'sd1219, 12'sd-1698, 11'sd751}},
{{11'sd849, 11'sd778, 12'sd1676}, {13'sd-2093, 10'sd343, 13'sd2481}, {12'sd-1503, 10'sd-350, 11'sd985}},
{{12'sd1152, 12'sd-1078, 13'sd-3092}, {13'sd-2632, 12'sd-1901, 11'sd705}, {11'sd518, 9'sd214, 12'sd-1905}},
{{12'sd-1375, 13'sd2361, 11'sd937}, {12'sd-1618, 12'sd1333, 6'sd26}, {9'sd-170, 11'sd-843, 11'sd514}},
{{12'sd1892, 10'sd295, 12'sd1286}, {9'sd186, 13'sd2193, 13'sd2320}, {12'sd-1219, 11'sd-746, 13'sd-2464}},
{{10'sd448, 8'sd118, 11'sd-525}, {10'sd-320, 13'sd-2972, 12'sd-1141}, {12'sd-1907, 9'sd229, 12'sd-1616}},
{{11'sd530, 12'sd1133, 12'sd1581}, {11'sd-990, 13'sd2704, 12'sd1118}, {13'sd2490, 10'sd432, 13'sd2069}},
{{13'sd2363, 13'sd2240, 11'sd573}, {13'sd3068, 13'sd-2229, 11'sd587}, {12'sd1280, 13'sd3089, 12'sd1183}},
{{11'sd518, 11'sd-741, 11'sd550}, {12'sd-1816, 13'sd2735, 12'sd-1934}, {7'sd59, 9'sd155, 12'sd1491}},
{{11'sd-781, 12'sd-1710, 11'sd-914}, {9'sd245, 8'sd-98, 13'sd3304}, {13'sd2576, 10'sd-335, 12'sd-1190}},
{{10'sd-444, 12'sd-1959, 13'sd-2329}, {13'sd-3013, 12'sd2042, 12'sd-1780}, {8'sd79, 13'sd-2272, 12'sd1670}},
{{13'sd2516, 12'sd1162, 13'sd-3072}, {11'sd682, 12'sd-1367, 13'sd-2650}, {13'sd2167, 12'sd-1862, 10'sd465}},
{{12'sd1886, 10'sd430, 13'sd3343}, {11'sd-911, 12'sd1944, 13'sd3303}, {13'sd3228, 11'sd788, 12'sd1367}},
{{11'sd743, 12'sd-1894, 10'sd286}, {10'sd-306, 12'sd1066, 12'sd1420}, {7'sd51, 13'sd2287, 13'sd2599}},
{{12'sd1166, 9'sd219, 12'sd-1680}, {13'sd2725, 13'sd3206, 12'sd-1406}, {12'sd1793, 9'sd-186, 12'sd1588}},
{{11'sd-959, 11'sd832, 10'sd-441}, {13'sd-2379, 11'sd-980, 10'sd488}, {12'sd-1781, 13'sd-2735, 8'sd117}},
{{12'sd1766, 11'sd-979, 10'sd-282}, {12'sd1979, 12'sd1575, 12'sd1110}, {13'sd-2353, 6'sd24, 12'sd1091}},
{{12'sd-2001, 11'sd-957, 13'sd-2173}, {13'sd-2220, 12'sd-1617, 13'sd2640}, {11'sd880, 12'sd1489, 13'sd2729}},
{{12'sd-2029, 13'sd2352, 11'sd-917}, {12'sd-1707, 7'sd35, 12'sd1579}, {8'sd107, 9'sd149, 8'sd-121}},
{{13'sd-2270, 10'sd-333, 12'sd1229}, {13'sd-2896, 12'sd-1058, 11'sd728}, {11'sd656, 13'sd-3801, 3'sd3}},
{{13'sd-2988, 13'sd-2195, 10'sd-511}, {13'sd-2277, 10'sd-299, 12'sd-1659}, {12'sd-1816, 11'sd-744, 6'sd-26}},
{{10'sd312, 9'sd-140, 12'sd1204}, {12'sd1532, 11'sd522, 11'sd686}, {12'sd1255, 12'sd1781, 12'sd1212}},
{{11'sd922, 8'sd-65, 12'sd-1727}, {13'sd2651, 6'sd-19, 12'sd-1904}, {11'sd776, 13'sd2376, 12'sd1294}},
{{12'sd-1423, 13'sd-2085, 13'sd2273}, {12'sd1400, 12'sd-1700, 13'sd-2451}, {11'sd-603, 13'sd-2138, 13'sd-2090}},
{{13'sd-2334, 13'sd-2226, 13'sd2172}, {12'sd-1924, 11'sd790, 13'sd2222}, {13'sd-2566, 12'sd1549, 9'sd-172}},
{{9'sd193, 12'sd1848, 13'sd2070}, {13'sd2080, 12'sd-1994, 12'sd-1238}, {9'sd242, 11'sd939, 12'sd-1972}},
{{13'sd-2935, 11'sd517, 13'sd-2133}, {12'sd2044, 11'sd-987, 13'sd-2116}, {12'sd1148, 11'sd-584, 12'sd-1053}},
{{12'sd-1808, 13'sd2681, 7'sd36}, {12'sd-1773, 12'sd-1363, 8'sd-98}, {13'sd-2872, 12'sd-1935, 12'sd-1373}},
{{13'sd-2187, 13'sd2379, 13'sd-2682}, {11'sd-665, 13'sd-2776, 13'sd-2281}, {12'sd-1939, 13'sd2425, 13'sd-2585}},
{{12'sd1767, 11'sd753, 13'sd-3183}, {12'sd-1775, 13'sd-2265, 12'sd1199}, {13'sd2245, 13'sd3266, 12'sd1809}},
{{11'sd985, 9'sd251, 13'sd-2366}, {12'sd-1815, 13'sd-2320, 10'sd266}, {11'sd530, 12'sd1912, 13'sd2179}},
{{8'sd71, 8'sd-120, 12'sd1295}, {11'sd-531, 12'sd-2042, 13'sd-2597}, {12'sd1780, 11'sd578, 13'sd2137}},
{{12'sd-1051, 13'sd2405, 11'sd591}, {13'sd-2187, 10'sd-298, 13'sd2136}, {12'sd1926, 13'sd2155, 13'sd-2273}},
{{12'sd-1356, 13'sd2100, 12'sd-1531}, {11'sd632, 10'sd-402, 12'sd-1251}, {12'sd-1609, 10'sd-487, 13'sd2554}},
{{13'sd2231, 11'sd960, 12'sd1144}, {12'sd1063, 12'sd-1871, 11'sd571}, {12'sd1625, 11'sd746, 11'sd-787}},
{{12'sd1181, 9'sd180, 13'sd-2152}, {13'sd2439, 13'sd2083, 12'sd-1415}, {11'sd1004, 12'sd1988, 12'sd1174}},
{{10'sd300, 9'sd153, 11'sd-736}, {13'sd2800, 11'sd749, 13'sd2200}, {10'sd-390, 12'sd-1222, 13'sd-3219}},
{{13'sd2417, 12'sd-1506, 11'sd-597}, {12'sd1891, 12'sd-1700, 13'sd-2472}, {10'sd431, 12'sd-1264, 12'sd-1966}},
{{11'sd-916, 13'sd-2628, 12'sd-1876}, {12'sd1366, 10'sd-321, 11'sd-699}, {13'sd-2138, 13'sd2176, 13'sd-2225}},
{{12'sd1767, 11'sd-561, 11'sd-931}, {12'sd-1182, 11'sd-910, 13'sd2734}, {11'sd-654, 12'sd-1216, 12'sd1928}},
{{12'sd-1360, 12'sd1115, 12'sd-1393}, {12'sd-1918, 11'sd618, 12'sd1213}, {8'sd-99, 13'sd-2295, 13'sd2690}},
{{11'sd-647, 11'sd855, 13'sd-2707}, {11'sd-658, 9'sd-134, 12'sd1402}, {10'sd355, 12'sd1296, 11'sd-527}},
{{10'sd339, 12'sd1039, 12'sd-1196}, {9'sd244, 13'sd-2285, 12'sd-1054}, {11'sd-737, 11'sd-573, 6'sd25}}},
{
{{10'sd262, 11'sd977, 12'sd-1833}, {13'sd-2396, 13'sd-2573, 11'sd886}, {13'sd-2634, 13'sd-2200, 9'sd-188}},
{{13'sd2675, 12'sd-1381, 12'sd-1894}, {12'sd-1170, 13'sd-2341, 12'sd1878}, {12'sd-1210, 12'sd-1488, 11'sd669}},
{{12'sd-1347, 12'sd1634, 11'sd-796}, {11'sd905, 12'sd1486, 12'sd-1484}, {5'sd11, 9'sd-251, 11'sd-993}},
{{13'sd-2269, 9'sd-145, 13'sd-2400}, {13'sd-2935, 13'sd-2982, 10'sd440}, {10'sd361, 11'sd-546, 12'sd-2044}},
{{11'sd591, 13'sd2938, 12'sd-1261}, {10'sd480, 12'sd-1444, 12'sd-1447}, {13'sd2675, 12'sd1258, 10'sd457}},
{{13'sd2547, 12'sd1250, 12'sd1309}, {13'sd2678, 12'sd-1979, 12'sd-1993}, {13'sd2090, 12'sd1080, 12'sd1579}},
{{13'sd2969, 12'sd1127, 12'sd-1324}, {12'sd-1067, 12'sd-1313, 9'sd-245}, {11'sd-659, 12'sd-1162, 6'sd-18}},
{{11'sd-958, 12'sd1874, 11'sd792}, {10'sd-450, 13'sd2592, 10'sd-433}, {13'sd-2525, 12'sd1148, 12'sd1857}},
{{10'sd333, 9'sd149, 11'sd-1008}, {11'sd-525, 11'sd729, 11'sd861}, {13'sd2061, 9'sd139, 8'sd-81}},
{{11'sd-717, 10'sd385, 10'sd305}, {12'sd-1509, 9'sd158, 11'sd964}, {12'sd1827, 11'sd-644, 12'sd1274}},
{{13'sd-2890, 9'sd-152, 13'sd2141}, {10'sd373, 11'sd-657, 11'sd927}, {13'sd2525, 12'sd1450, 10'sd-462}},
{{12'sd1287, 12'sd1757, 13'sd2218}, {6'sd21, 10'sd-415, 12'sd1749}, {12'sd-1258, 13'sd-2567, 12'sd1568}},
{{13'sd3689, 10'sd-351, 7'sd38}, {12'sd1686, 13'sd-3382, 12'sd-1753}, {11'sd-652, 13'sd-3121, 14'sd-4358}},
{{13'sd3053, 12'sd1056, 11'sd574}, {12'sd1482, 12'sd1403, 13'sd-2660}, {12'sd-1448, 11'sd565, 13'sd2333}},
{{13'sd-2426, 7'sd-39, 12'sd-1024}, {12'sd-1531, 13'sd2201, 11'sd605}, {11'sd-619, 12'sd1024, 12'sd-1255}},
{{10'sd-290, 11'sd687, 12'sd1291}, {11'sd-850, 11'sd763, 13'sd-2270}, {12'sd1324, 12'sd-1993, 4'sd7}},
{{13'sd-2234, 13'sd3056, 12'sd1161}, {12'sd-1063, 12'sd1035, 11'sd982}, {12'sd1169, 12'sd-1563, 11'sd740}},
{{13'sd-2862, 9'sd-232, 13'sd-2722}, {11'sd-917, 12'sd1579, 10'sd352}, {12'sd-1520, 13'sd2745, 11'sd-587}},
{{10'sd379, 13'sd-2156, 13'sd2559}, {12'sd2021, 13'sd2585, 12'sd1267}, {12'sd1110, 12'sd-2043, 11'sd-873}},
{{12'sd1418, 13'sd-2469, 13'sd2909}, {12'sd2036, 12'sd-1060, 13'sd2254}, {13'sd3031, 13'sd2331, 11'sd-842}},
{{12'sd1622, 12'sd1802, 9'sd-211}, {12'sd-2033, 12'sd-1620, 11'sd533}, {8'sd-68, 11'sd897, 13'sd2553}},
{{11'sd852, 9'sd-215, 12'sd1966}, {13'sd-2159, 13'sd-2115, 13'sd-2082}, {10'sd271, 11'sd-928, 12'sd-1321}},
{{13'sd2722, 13'sd-2048, 7'sd-56}, {12'sd1659, 12'sd1962, 10'sd410}, {13'sd-2691, 10'sd-482, 12'sd1887}},
{{12'sd-1965, 12'sd-1745, 11'sd-908}, {11'sd-916, 10'sd484, 11'sd-833}, {12'sd-1134, 11'sd-779, 9'sd-187}},
{{10'sd-328, 7'sd-44, 11'sd-845}, {12'sd-1667, 12'sd1721, 13'sd2116}, {11'sd-1009, 9'sd-237, 13'sd3008}},
{{11'sd993, 12'sd1944, 11'sd-944}, {11'sd-652, 13'sd2501, 12'sd-1709}, {12'sd-1494, 8'sd-78, 12'sd1492}},
{{13'sd-2821, 13'sd-2679, 13'sd-2462}, {13'sd-2581, 10'sd-410, 10'sd473}, {12'sd1747, 8'sd109, 11'sd964}},
{{11'sd855, 12'sd1026, 11'sd-598}, {12'sd1593, 12'sd1634, 12'sd1175}, {10'sd-345, 11'sd1002, 13'sd-2379}},
{{13'sd2475, 10'sd403, 11'sd-688}, {13'sd-2401, 13'sd-2584, 11'sd-812}, {13'sd-2946, 12'sd-1482, 13'sd2667}},
{{12'sd-1987, 12'sd-1794, 12'sd1804}, {12'sd-1261, 12'sd1609, 13'sd2147}, {10'sd-320, 12'sd1183, 11'sd-907}},
{{13'sd-2891, 13'sd2592, 11'sd-854}, {13'sd-2248, 13'sd3206, 12'sd1958}, {8'sd118, 12'sd1712, 13'sd3186}},
{{13'sd2423, 12'sd1834, 11'sd776}, {12'sd-1466, 12'sd1543, 10'sd338}, {12'sd1335, 12'sd-1609, 10'sd-481}},
{{9'sd201, 13'sd-2661, 13'sd-2074}, {13'sd-3500, 13'sd-2904, 13'sd-2371}, {13'sd-3834, 12'sd-1778, 13'sd-2238}},
{{13'sd3425, 11'sd598, 8'sd111}, {12'sd1752, 12'sd1669, 12'sd-1893}, {6'sd-24, 13'sd2058, 13'sd2756}},
{{12'sd1045, 11'sd-612, 13'sd2109}, {13'sd2373, 11'sd-872, 11'sd-904}, {8'sd-121, 7'sd51, 12'sd1634}},
{{11'sd813, 11'sd-693, 12'sd1984}, {11'sd-965, 13'sd2614, 9'sd-205}, {12'sd1372, 12'sd1807, 13'sd2910}},
{{10'sd-411, 12'sd1995, 13'sd2674}, {11'sd-828, 10'sd315, 12'sd1944}, {13'sd2564, 13'sd2334, 12'sd-1035}},
{{13'sd2115, 12'sd-1162, 11'sd715}, {11'sd-623, 12'sd-1187, 10'sd-478}, {11'sd-552, 12'sd-1892, 12'sd1385}},
{{12'sd-1276, 12'sd-1942, 12'sd1297}, {13'sd2479, 7'sd34, 13'sd-2990}, {11'sd946, 11'sd752, 13'sd-2324}},
{{13'sd-2684, 6'sd-25, 11'sd-528}, {12'sd-1549, 11'sd-966, 13'sd2242}, {12'sd1796, 10'sd-360, 13'sd2336}},
{{13'sd-2503, 12'sd-1158, 12'sd-1296}, {9'sd-155, 12'sd-1760, 9'sd203}, {12'sd1927, 13'sd2998, 12'sd1584}},
{{13'sd2835, 10'sd-399, 11'sd808}, {10'sd-359, 13'sd2503, 12'sd1515}, {12'sd-1705, 12'sd1996, 12'sd1952}},
{{11'sd926, 11'sd-729, 11'sd-774}, {10'sd-390, 11'sd641, 13'sd-2881}, {13'sd2259, 11'sd845, 11'sd-850}},
{{11'sd595, 12'sd-1268, 7'sd-46}, {13'sd-2424, 13'sd-2114, 12'sd1945}, {9'sd-255, 13'sd2568, 10'sd430}},
{{12'sd1263, 9'sd255, 13'sd2224}, {13'sd-2085, 12'sd-1589, 12'sd1101}, {13'sd2138, 12'sd-1050, 8'sd-73}},
{{13'sd2094, 12'sd1953, 12'sd1494}, {8'sd-117, 11'sd-597, 13'sd-2137}, {10'sd-367, 6'sd-29, 12'sd1451}},
{{8'sd-115, 12'sd-1960, 13'sd-2318}, {12'sd1467, 12'sd-1201, 12'sd1662}, {13'sd2476, 10'sd-271, 8'sd-68}},
{{12'sd1440, 13'sd3325, 11'sd-819}, {11'sd563, 12'sd-1964, 12'sd2015}, {13'sd2472, 12'sd1442, 12'sd-1316}},
{{12'sd-1832, 11'sd-582, 10'sd364}, {13'sd-3201, 12'sd2009, 12'sd-1346}, {10'sd333, 11'sd717, 12'sd-1156}},
{{10'sd-429, 12'sd-1449, 12'sd1329}, {13'sd-2644, 10'sd-333, 12'sd1287}, {13'sd2254, 13'sd2591, 11'sd-565}},
{{12'sd1899, 12'sd1466, 12'sd-1626}, {12'sd-1159, 11'sd683, 12'sd1757}, {12'sd-1621, 13'sd-2057, 13'sd-3404}},
{{11'sd-617, 13'sd-2994, 13'sd2166}, {12'sd1572, 12'sd1251, 12'sd-1252}, {12'sd1425, 13'sd-2157, 11'sd-525}},
{{9'sd154, 13'sd-2438, 12'sd1818}, {11'sd-564, 11'sd793, 11'sd-953}, {12'sd-1717, 10'sd377, 9'sd-249}},
{{12'sd-1287, 11'sd757, 11'sd-923}, {11'sd-659, 12'sd-1384, 12'sd1860}, {13'sd-2741, 12'sd1535, 13'sd-2688}},
{{12'sd1706, 12'sd1242, 11'sd569}, {13'sd-2419, 12'sd-1347, 11'sd-985}, {12'sd-1461, 9'sd160, 13'sd-3108}},
{{12'sd-1690, 13'sd2546, 7'sd55}, {9'sd189, 11'sd-892, 12'sd1848}, {10'sd-426, 11'sd-704, 11'sd-766}},
{{9'sd144, 12'sd1517, 12'sd1240}, {8'sd86, 12'sd-1663, 12'sd-2010}, {7'sd-33, 11'sd787, 11'sd-703}},
{{13'sd3050, 11'sd642, 11'sd896}, {13'sd2914, 12'sd1427, 13'sd2284}, {8'sd-102, 10'sd-384, 13'sd-2098}},
{{13'sd2128, 7'sd60, 12'sd-1381}, {10'sd342, 13'sd-2341, 12'sd1416}, {12'sd-1941, 11'sd642, 8'sd94}},
{{13'sd3662, 13'sd3249, 11'sd745}, {12'sd-1498, 13'sd-2732, 12'sd-1187}, {13'sd2410, 11'sd593, 12'sd-1926}},
{{13'sd-2426, 11'sd-553, 12'sd-1460}, {10'sd349, 11'sd-716, 11'sd-879}, {11'sd-704, 9'sd-155, 12'sd1334}},
{{12'sd-1558, 12'sd-1872, 13'sd-2701}, {13'sd-2180, 13'sd-2220, 13'sd2675}, {11'sd-931, 12'sd1933, 8'sd127}},
{{9'sd215, 8'sd-111, 12'sd-1330}, {12'sd-1818, 13'sd2277, 12'sd-1409}, {13'sd-2652, 13'sd-2488, 7'sd-33}},
{{11'sd-648, 11'sd-716, 12'sd1447}, {11'sd-844, 11'sd836, 11'sd677}, {13'sd2386, 11'sd974, 11'sd728}}},
{
{{11'sd-946, 12'sd1649, 12'sd1502}, {4'sd7, 10'sd402, 11'sd-571}, {12'sd1400, 9'sd212, 8'sd116}},
{{12'sd1195, 10'sd-441, 11'sd-870}, {13'sd2337, 12'sd1184, 12'sd1991}, {8'sd93, 12'sd-1877, 12'sd-1580}},
{{11'sd-642, 13'sd-2904, 10'sd-500}, {6'sd-28, 13'sd2190, 12'sd-1240}, {13'sd-3589, 13'sd-2532, 13'sd2347}},
{{11'sd-951, 12'sd-1069, 10'sd-313}, {8'sd-76, 10'sd268, 10'sd294}, {5'sd-10, 10'sd-313, 11'sd-820}},
{{12'sd1394, 13'sd2289, 12'sd-1404}, {11'sd-843, 11'sd907, 11'sd670}, {12'sd1045, 10'sd494, 11'sd-910}},
{{12'sd-1891, 11'sd-976, 10'sd320}, {11'sd621, 13'sd-2049, 13'sd2630}, {10'sd315, 10'sd-468, 13'sd2669}},
{{11'sd1017, 11'sd-877, 11'sd989}, {13'sd2754, 9'sd-215, 12'sd1531}, {14'sd4504, 12'sd1382, 13'sd2206}},
{{11'sd-633, 11'sd-942, 13'sd3108}, {13'sd2111, 12'sd1469, 13'sd3417}, {13'sd-2104, 12'sd1589, 11'sd-603}},
{{11'sd-1007, 12'sd1052, 12'sd-1647}, {10'sd-350, 13'sd2435, 13'sd-2429}, {8'sd-114, 13'sd-2305, 13'sd-2055}},
{{12'sd-1429, 13'sd2111, 12'sd-1609}, {10'sd-318, 11'sd676, 12'sd1458}, {10'sd-287, 10'sd257, 10'sd-306}},
{{13'sd-2886, 11'sd517, 12'sd1330}, {13'sd2477, 10'sd292, 13'sd2674}, {8'sd-117, 11'sd830, 12'sd1945}},
{{13'sd-2494, 13'sd-2251, 11'sd967}, {12'sd-1263, 12'sd1791, 11'sd-628}, {9'sd-223, 13'sd2074, 12'sd1370}},
{{11'sd-630, 13'sd-2106, 14'sd-7021}, {13'sd2367, 11'sd1015, 12'sd-1475}, {12'sd1545, 12'sd-1554, 12'sd1088}},
{{11'sd949, 11'sd813, 13'sd2285}, {9'sd131, 13'sd-2100, 11'sd812}, {12'sd1718, 13'sd2125, 13'sd-2061}},
{{12'sd1597, 11'sd-612, 12'sd-1769}, {12'sd-1597, 13'sd2582, 13'sd-3140}, {13'sd2119, 12'sd-1799, 13'sd-3022}},
{{13'sd2556, 13'sd2285, 13'sd2244}, {11'sd-854, 13'sd-2226, 9'sd141}, {13'sd2121, 11'sd-813, 13'sd3164}},
{{12'sd-1718, 11'sd1007, 11'sd992}, {12'sd1523, 12'sd-1109, 12'sd1843}, {8'sd-127, 11'sd-919, 12'sd-1964}},
{{7'sd-36, 12'sd1949, 12'sd-1486}, {7'sd-61, 13'sd2531, 13'sd-2338}, {13'sd-2320, 11'sd619, 12'sd-2017}},
{{13'sd-2455, 13'sd-3072, 8'sd107}, {12'sd-1952, 13'sd-2099, 13'sd-3025}, {12'sd-1428, 11'sd-840, 13'sd2060}},
{{12'sd1542, 12'sd-1467, 12'sd-1949}, {11'sd912, 12'sd-1062, 10'sd-498}, {12'sd2013, 13'sd2330, 11'sd-661}},
{{10'sd269, 13'sd3538, 12'sd1689}, {13'sd2841, 11'sd-742, 13'sd2998}, {9'sd-187, 11'sd717, 13'sd2208}},
{{13'sd-2406, 12'sd-1699, 13'sd-3667}, {13'sd-2149, 10'sd334, 11'sd-844}, {11'sd-613, 12'sd-1097, 13'sd2760}},
{{8'sd-103, 12'sd-1304, 12'sd-1123}, {11'sd923, 11'sd872, 13'sd-2369}, {12'sd-1439, 13'sd-2480, 12'sd-1449}},
{{10'sd289, 12'sd1302, 11'sd571}, {12'sd-1686, 12'sd1877, 13'sd-2776}, {11'sd-664, 12'sd-1142, 13'sd-2298}},
{{13'sd2059, 13'sd-2670, 13'sd2368}, {12'sd1490, 13'sd-2277, 12'sd-1038}, {13'sd2900, 13'sd2572, 13'sd2612}},
{{13'sd2665, 13'sd2305, 8'sd79}, {8'sd-82, 12'sd1320, 11'sd624}, {12'sd1959, 13'sd2887, 12'sd1581}},
{{12'sd1926, 12'sd-1992, 12'sd1421}, {12'sd1227, 12'sd-1388, 12'sd-1863}, {13'sd-2212, 13'sd-2590, 12'sd1626}},
{{13'sd2273, 9'sd-194, 11'sd-518}, {12'sd1897, 12'sd-1704, 9'sd-133}, {8'sd-124, 10'sd-278, 12'sd1408}},
{{12'sd-1916, 11'sd-655, 12'sd-1398}, {12'sd1841, 12'sd-1794, 12'sd1354}, {12'sd-1584, 12'sd1788, 12'sd1394}},
{{13'sd-2055, 12'sd-1463, 12'sd1778}, {13'sd2820, 8'sd-119, 13'sd-2366}, {13'sd-2364, 12'sd1390, 12'sd-1363}},
{{11'sd-751, 11'sd-978, 10'sd-425}, {12'sd1417, 13'sd2759, 12'sd-1350}, {13'sd2867, 13'sd2746, 13'sd2954}},
{{12'sd1318, 13'sd2863, 11'sd972}, {11'sd-632, 11'sd628, 12'sd1553}, {12'sd1081, 12'sd1713, 12'sd-1335}},
{{11'sd-888, 10'sd398, 11'sd928}, {11'sd-786, 11'sd-550, 12'sd1401}, {11'sd-534, 8'sd115, 13'sd3033}},
{{13'sd2233, 11'sd-993, 13'sd3437}, {9'sd-224, 12'sd1187, 11'sd899}, {11'sd785, 11'sd-840, 12'sd-1144}},
{{12'sd1183, 11'sd-946, 12'sd1550}, {5'sd11, 12'sd1065, 13'sd2057}, {11'sd975, 13'sd-2659, 13'sd2099}},
{{13'sd-2845, 12'sd1472, 10'sd272}, {12'sd1333, 11'sd-925, 13'sd-2054}, {12'sd-1466, 12'sd-2019, 12'sd1385}},
{{12'sd-1590, 12'sd-2009, 11'sd590}, {13'sd-2399, 11'sd993, 13'sd2134}, {12'sd-1710, 11'sd561, 9'sd176}},
{{12'sd-1754, 13'sd-2141, 11'sd740}, {12'sd-1837, 12'sd-1957, 12'sd-1570}, {13'sd2344, 13'sd-2311, 12'sd-1583}},
{{13'sd3842, 13'sd2066, 12'sd1844}, {10'sd407, 9'sd-186, 12'sd1604}, {12'sd-1758, 13'sd-2807, 12'sd1805}},
{{12'sd-1812, 13'sd2264, 12'sd1555}, {13'sd-2272, 13'sd2327, 12'sd1688}, {9'sd-236, 13'sd2102, 13'sd-2211}},
{{11'sd-641, 11'sd658, 10'sd485}, {13'sd-4043, 8'sd-117, 11'sd-627}, {8'sd-82, 13'sd2954, 8'sd79}},
{{10'sd-417, 13'sd-2939, 13'sd-3431}, {9'sd253, 11'sd-733, 11'sd-780}, {11'sd658, 4'sd6, 12'sd1461}},
{{11'sd-822, 12'sd1889, 11'sd-647}, {12'sd2035, 10'sd-456, 11'sd-944}, {13'sd-2162, 11'sd907, 13'sd2369}},
{{13'sd-2520, 13'sd-2595, 11'sd-642}, {13'sd2095, 11'sd667, 11'sd-552}, {10'sd480, 13'sd-2888, 13'sd-2265}},
{{11'sd-823, 11'sd-931, 4'sd6}, {12'sd-1365, 12'sd1670, 12'sd-1271}, {12'sd-1431, 12'sd1779, 13'sd2605}},
{{13'sd-2124, 10'sd-491, 8'sd-96}, {12'sd-1904, 13'sd-2276, 13'sd-2339}, {13'sd-2710, 10'sd-507, 11'sd590}},
{{10'sd302, 12'sd1061, 13'sd-2091}, {13'sd-2564, 13'sd2147, 13'sd2452}, {12'sd1400, 13'sd-2883, 13'sd2384}},
{{12'sd1169, 13'sd-3147, 13'sd-3046}, {12'sd1891, 10'sd-290, 12'sd-1133}, {12'sd-1909, 13'sd-3462, 13'sd-3635}},
{{13'sd2450, 12'sd-1577, 13'sd2500}, {12'sd-2006, 12'sd1238, 12'sd2030}, {12'sd-1552, 13'sd2626, 11'sd-603}},
{{13'sd-3099, 8'sd-116, 10'sd-458}, {14'sd-4174, 9'sd205, 13'sd-2641}, {10'sd333, 11'sd979, 13'sd-2517}},
{{12'sd-1155, 8'sd-89, 12'sd-1926}, {12'sd1602, 13'sd-3186, 9'sd227}, {9'sd187, 13'sd-2717, 11'sd865}},
{{12'sd-1815, 10'sd403, 10'sd-488}, {10'sd417, 12'sd-1602, 11'sd768}, {12'sd-1593, 13'sd-2400, 13'sd-2372}},
{{12'sd1520, 12'sd1720, 12'sd-1564}, {12'sd-1190, 12'sd1075, 10'sd332}, {12'sd1795, 11'sd-751, 11'sd-773}},
{{11'sd732, 11'sd-836, 9'sd-226}, {11'sd850, 13'sd2497, 13'sd2769}, {13'sd2550, 12'sd1951, 13'sd2506}},
{{11'sd-904, 12'sd-1260, 8'sd81}, {12'sd1038, 12'sd1617, 13'sd3040}, {12'sd-1542, 11'sd977, 13'sd2657}},
{{12'sd1070, 11'sd714, 12'sd1172}, {13'sd2171, 11'sd-981, 12'sd-1860}, {12'sd-1520, 10'sd-281, 12'sd1342}},
{{12'sd1426, 13'sd2472, 12'sd1116}, {12'sd-1220, 9'sd-233, 11'sd882}, {12'sd-1325, 10'sd-435, 12'sd-1256}},
{{12'sd-1422, 11'sd788, 13'sd-3188}, {13'sd2101, 14'sd4103, 11'sd830}, {12'sd1173, 13'sd2469, 13'sd-3565}},
{{10'sd-264, 11'sd1008, 13'sd2060}, {13'sd2160, 13'sd-3238, 11'sd-619}, {11'sd829, 11'sd791, 12'sd1364}},
{{13'sd2388, 12'sd-1149, 11'sd-923}, {13'sd3785, 13'sd-2637, 13'sd3422}, {12'sd1837, 11'sd776, 12'sd1724}},
{{11'sd726, 12'sd-1851, 13'sd-2755}, {10'sd-317, 12'sd1029, 11'sd-839}, {11'sd-542, 13'sd-2603, 12'sd-1215}},
{{12'sd-1962, 11'sd1003, 12'sd-1375}, {12'sd2034, 12'sd-1318, 11'sd-948}, {11'sd-875, 12'sd1968, 11'sd-523}},
{{12'sd2017, 11'sd-776, 12'sd-1564}, {11'sd638, 12'sd-1201, 12'sd1906}, {12'sd-1675, 10'sd423, 12'sd1211}},
{{12'sd1980, 12'sd1944, 11'sd671}, {12'sd1977, 12'sd-1250, 13'sd-2324}, {12'sd-1289, 10'sd414, 13'sd-2750}}},
{
{{12'sd-1618, 11'sd-699, 12'sd1171}, {12'sd1465, 8'sd-88, 13'sd-2387}, {12'sd-1907, 13'sd-2601, 12'sd-1084}},
{{13'sd2202, 12'sd-1758, 12'sd1639}, {11'sd-580, 12'sd1490, 7'sd47}, {12'sd1236, 11'sd-975, 12'sd1176}},
{{11'sd936, 12'sd-1983, 13'sd-2858}, {12'sd-1443, 13'sd3335, 11'sd-562}, {13'sd-3158, 8'sd-69, 11'sd-922}},
{{13'sd2383, 11'sd628, 12'sd1346}, {8'sd105, 12'sd-1198, 13'sd-2268}, {14'sd-4613, 12'sd1073, 13'sd-3015}},
{{12'sd-1972, 12'sd1759, 13'sd2441}, {11'sd-855, 12'sd-1429, 13'sd-2172}, {11'sd-701, 10'sd418, 13'sd-2211}},
{{12'sd1276, 11'sd719, 13'sd2133}, {13'sd2359, 12'sd1610, 13'sd-2282}, {12'sd-1620, 13'sd-2579, 13'sd-2541}},
{{12'sd1182, 12'sd-1704, 13'sd-2505}, {12'sd-1966, 12'sd-1878, 10'sd-478}, {13'sd2100, 13'sd2321, 13'sd3931}},
{{11'sd970, 12'sd-1500, 10'sd493}, {13'sd2652, 10'sd272, 10'sd-359}, {13'sd-3272, 13'sd2731, 13'sd-2641}},
{{10'sd450, 13'sd2070, 13'sd2417}, {11'sd724, 13'sd3231, 10'sd-319}, {13'sd-2218, 13'sd2048, 9'sd-182}},
{{13'sd-2505, 11'sd-901, 12'sd-1882}, {13'sd2084, 11'sd759, 11'sd-520}, {12'sd1687, 12'sd1530, 8'sd-90}},
{{10'sd-295, 12'sd-1104, 13'sd2379}, {12'sd1089, 12'sd-1361, 12'sd-1740}, {12'sd-1056, 11'sd-622, 13'sd2603}},
{{11'sd-547, 13'sd-2921, 10'sd-396}, {12'sd1433, 10'sd413, 11'sd884}, {11'sd1020, 11'sd-624, 10'sd312}},
{{14'sd-4799, 10'sd-317, 13'sd-3520}, {13'sd3510, 11'sd-1019, 11'sd912}, {8'sd102, 11'sd698, 12'sd1906}},
{{12'sd-1385, 12'sd-1904, 12'sd1731}, {10'sd418, 12'sd1910, 12'sd1971}, {9'sd-221, 12'sd1466, 11'sd893}},
{{12'sd1504, 13'sd-2145, 12'sd-1580}, {13'sd2497, 12'sd-1492, 10'sd-488}, {13'sd2198, 12'sd-1383, 5'sd-8}},
{{13'sd2532, 12'sd-1614, 13'sd2613}, {13'sd2710, 11'sd-699, 13'sd2259}, {12'sd1319, 12'sd-1987, 12'sd-1452}},
{{13'sd2494, 12'sd1213, 7'sd-33}, {12'sd1722, 9'sd229, 9'sd-158}, {11'sd-1021, 11'sd-825, 7'sd43}},
{{12'sd1418, 13'sd3089, 8'sd123}, {11'sd814, 13'sd2810, 12'sd1222}, {9'sd228, 11'sd614, 12'sd-1254}},
{{13'sd-2423, 12'sd1600, 11'sd960}, {12'sd-1507, 10'sd-380, 13'sd2120}, {11'sd888, 12'sd2029, 12'sd-1559}},
{{12'sd1403, 13'sd-2378, 13'sd-2054}, {13'sd3174, 12'sd-1024, 7'sd52}, {11'sd516, 8'sd-76, 9'sd-177}},
{{12'sd1962, 13'sd3055, 11'sd654}, {13'sd2192, 11'sd743, 12'sd-1467}, {12'sd-1467, 12'sd1796, 12'sd-1480}},
{{13'sd-2626, 11'sd933, 13'sd-3134}, {10'sd287, 12'sd1190, 11'sd774}, {12'sd1335, 13'sd-2504, 13'sd3302}},
{{12'sd1463, 11'sd581, 10'sd434}, {13'sd-2097, 13'sd2583, 12'sd1109}, {9'sd240, 11'sd-569, 13'sd-3622}},
{{13'sd2333, 12'sd-1374, 12'sd-1983}, {9'sd-226, 10'sd-379, 11'sd978}, {11'sd989, 11'sd537, 13'sd-3210}},
{{11'sd-834, 12'sd-1734, 11'sd585}, {11'sd-596, 13'sd-2238, 12'sd-1326}, {12'sd1205, 11'sd739, 10'sd-433}},
{{11'sd552, 13'sd-2067, 8'sd124}, {13'sd2864, 13'sd2775, 12'sd1587}, {11'sd633, 12'sd1037, 9'sd221}},
{{12'sd1647, 12'sd-1677, 12'sd1778}, {13'sd2260, 10'sd-478, 11'sd761}, {12'sd-1447, 12'sd-1419, 9'sd-250}},
{{12'sd1033, 11'sd955, 10'sd365}, {11'sd710, 11'sd-550, 11'sd-821}, {10'sd266, 12'sd-1688, 12'sd1977}},
{{12'sd1740, 13'sd-2224, 12'sd1857}, {12'sd1480, 11'sd603, 12'sd-1077}, {11'sd-1000, 12'sd1331, 13'sd-2170}},
{{10'sd-319, 12'sd1281, 13'sd2732}, {11'sd-943, 13'sd-2127, 12'sd-1231}, {10'sd284, 13'sd-2365, 12'sd-1612}},
{{11'sd-869, 13'sd3893, 11'sd936}, {13'sd2184, 12'sd1632, 7'sd-45}, {14'sd4906, 14'sd5666, 14'sd6310}},
{{13'sd2681, 13'sd2841, 11'sd-862}, {12'sd-1294, 13'sd2250, 5'sd9}, {10'sd-290, 11'sd-1023, 12'sd-1362}},
{{8'sd80, 12'sd-1800, 12'sd-1576}, {11'sd-828, 11'sd-851, 12'sd-1864}, {13'sd-3402, 12'sd1835, 13'sd2278}},
{{13'sd2283, 8'sd94, 13'sd2780}, {11'sd750, 12'sd-1295, 10'sd478}, {12'sd1667, 8'sd67, 12'sd-2030}},
{{11'sd-972, 11'sd-875, 13'sd2104}, {12'sd-1551, 13'sd2125, 10'sd-425}, {13'sd2964, 11'sd-973, 12'sd1184}},
{{10'sd-481, 11'sd-787, 12'sd-1403}, {12'sd-1319, 13'sd2541, 12'sd-1165}, {12'sd-1296, 11'sd-829, 12'sd-1260}},
{{12'sd1723, 11'sd-634, 11'sd-570}, {11'sd-853, 12'sd-1244, 11'sd826}, {9'sd241, 11'sd768, 10'sd-270}},
{{12'sd-1574, 12'sd-1932, 12'sd-1298}, {13'sd2487, 13'sd2641, 9'sd167}, {11'sd-648, 12'sd1935, 10'sd418}},
{{11'sd-1022, 12'sd-1363, 12'sd-1273}, {11'sd-1003, 12'sd-1683, 12'sd1156}, {12'sd-1072, 13'sd2096, 12'sd1187}},
{{8'sd107, 11'sd628, 12'sd1632}, {8'sd122, 10'sd257, 13'sd-2773}, {12'sd-1355, 12'sd-1408, 12'sd1920}},
{{12'sd-1728, 12'sd-1489, 13'sd-2609}, {8'sd-92, 9'sd-234, 12'sd1083}, {9'sd197, 10'sd366, 12'sd1643}},
{{12'sd-1721, 10'sd417, 11'sd763}, {12'sd1352, 12'sd1056, 11'sd-673}, {11'sd-950, 13'sd2365, 11'sd-976}},
{{13'sd-2348, 13'sd2409, 12'sd1286}, {11'sd949, 11'sd764, 12'sd-1724}, {3'sd-2, 7'sd34, 13'sd2051}},
{{9'sd-131, 11'sd840, 12'sd-1705}, {12'sd1823, 12'sd-1704, 9'sd174}, {11'sd-549, 11'sd-655, 12'sd1080}},
{{12'sd1716, 12'sd-2030, 13'sd-3116}, {12'sd-1400, 12'sd-1827, 13'sd2535}, {13'sd2286, 12'sd-1238, 12'sd1415}},
{{13'sd2657, 13'sd-2556, 12'sd1590}, {13'sd2833, 9'sd-218, 12'sd1414}, {10'sd-392, 11'sd879, 12'sd1690}},
{{12'sd1381, 13'sd-2883, 12'sd-1476}, {12'sd1561, 13'sd2525, 12'sd1528}, {13'sd2795, 13'sd-2075, 9'sd193}},
{{13'sd-3162, 11'sd-1001, 12'sd1958}, {12'sd-1912, 13'sd2252, 11'sd-866}, {13'sd2402, 12'sd1657, 13'sd2186}},
{{12'sd-1500, 9'sd143, 13'sd2647}, {12'sd-1308, 12'sd-1646, 11'sd546}, {13'sd-2452, 11'sd-763, 13'sd-2893}},
{{12'sd-1903, 10'sd382, 13'sd2105}, {9'sd232, 10'sd-360, 12'sd1202}, {12'sd1697, 11'sd-856, 13'sd-2214}},
{{12'sd1340, 9'sd-246, 11'sd604}, {10'sd-270, 13'sd-2839, 10'sd473}, {13'sd-2240, 12'sd-1630, 11'sd-685}},
{{12'sd-1106, 8'sd113, 13'sd-2571}, {13'sd-2093, 11'sd723, 11'sd-523}, {12'sd-1392, 13'sd2179, 12'sd-1952}},
{{12'sd1638, 11'sd-857, 12'sd1838}, {13'sd2653, 10'sd-292, 11'sd779}, {10'sd-450, 12'sd-1163, 13'sd2123}},
{{12'sd1443, 11'sd933, 13'sd2391}, {11'sd-766, 11'sd563, 11'sd-1002}, {13'sd-2305, 11'sd-782, 12'sd-1896}},
{{12'sd1060, 12'sd-1209, 14'sd-4347}, {11'sd-805, 6'sd18, 12'sd-2040}, {12'sd-1556, 12'sd1463, 12'sd1938}},
{{12'sd-1874, 10'sd-362, 11'sd-871}, {13'sd3415, 12'sd2020, 12'sd-1165}, {12'sd1049, 13'sd-2773, 13'sd-2060}},
{{11'sd784, 11'sd943, 12'sd1049}, {13'sd-2443, 12'sd2008, 12'sd1142}, {12'sd-1572, 11'sd905, 10'sd359}},
{{11'sd782, 13'sd-2208, 12'sd-1937}, {12'sd1103, 13'sd2735, 14'sd4673}, {14'sd4161, 13'sd-2319, 12'sd-1028}},
{{12'sd-1563, 12'sd-1401, 11'sd-799}, {11'sd-797, 12'sd-1277, 12'sd1196}, {13'sd2135, 13'sd3164, 13'sd2634}},
{{10'sd-306, 13'sd-2876, 12'sd1470}, {11'sd835, 12'sd1051, 10'sd277}, {13'sd2186, 13'sd-2245, 13'sd2220}},
{{11'sd-537, 13'sd2131, 8'sd95}, {12'sd1563, 12'sd1334, 13'sd-2610}, {11'sd579, 13'sd2239, 9'sd132}},
{{12'sd-1865, 10'sd396, 11'sd719}, {13'sd-2177, 12'sd1074, 12'sd-1980}, {10'sd368, 12'sd-1220, 9'sd-178}},
{{12'sd2026, 12'sd1144, 13'sd-2114}, {12'sd-1805, 12'sd-1123, 13'sd2709}, {12'sd-1622, 12'sd1778, 13'sd-2577}},
{{13'sd-2389, 13'sd-2969, 10'sd-268}, {12'sd-1114, 12'sd1274, 8'sd109}, {10'sd-417, 12'sd-1978, 11'sd788}}},
{
{{2'sd-1, 12'sd-1653, 12'sd1921}, {12'sd-1383, 12'sd-1276, 12'sd1441}, {10'sd-426, 12'sd-1772, 10'sd494}},
{{12'sd1583, 13'sd-2502, 13'sd-2435}, {11'sd950, 12'sd-1325, 12'sd-1526}, {12'sd1435, 13'sd-2142, 12'sd-1942}},
{{6'sd-31, 11'sd-671, 13'sd-2611}, {13'sd-2167, 6'sd-30, 12'sd-1727}, {10'sd288, 12'sd-1669, 13'sd2421}},
{{6'sd-31, 12'sd-1896, 12'sd1533}, {11'sd-833, 10'sd-317, 11'sd514}, {13'sd2210, 10'sd282, 11'sd-882}},
{{9'sd129, 13'sd2491, 9'sd237}, {10'sd-498, 13'sd-2185, 12'sd-1233}, {10'sd419, 13'sd2077, 12'sd-1886}},
{{13'sd-2202, 9'sd190, 10'sd-500}, {12'sd-1104, 13'sd-2686, 10'sd-329}, {10'sd-287, 12'sd-1521, 10'sd342}},
{{11'sd-671, 4'sd-4, 12'sd2037}, {10'sd446, 13'sd-2356, 10'sd382}, {8'sd117, 11'sd758, 8'sd-127}},
{{13'sd-2369, 13'sd-2127, 12'sd-1664}, {13'sd2243, 13'sd-2379, 12'sd1872}, {10'sd490, 12'sd1456, 13'sd2664}},
{{13'sd-3004, 11'sd-840, 12'sd-1966}, {13'sd-3058, 13'sd-2302, 12'sd1655}, {13'sd-2886, 12'sd-1790, 13'sd2564}},
{{9'sd-206, 10'sd-327, 12'sd1825}, {12'sd-1507, 13'sd-2133, 6'sd17}, {11'sd572, 7'sd61, 12'sd-1770}},
{{10'sd359, 12'sd-1783, 11'sd788}, {12'sd-1504, 12'sd-1322, 12'sd1710}, {9'sd-136, 11'sd-621, 13'sd-2337}},
{{12'sd-1442, 12'sd-1080, 6'sd28}, {12'sd1078, 11'sd707, 13'sd2474}, {11'sd-1019, 10'sd392, 13'sd-2671}},
{{13'sd2434, 11'sd842, 11'sd-860}, {10'sd332, 11'sd551, 13'sd-2905}, {12'sd1481, 12'sd-1550, 12'sd1201}},
{{12'sd1134, 13'sd-2308, 13'sd2793}, {11'sd1023, 13'sd2180, 10'sd370}, {13'sd-2565, 12'sd-1593, 12'sd-1623}},
{{13'sd3264, 13'sd-2087, 12'sd-1401}, {13'sd2399, 12'sd1892, 12'sd1507}, {12'sd1089, 5'sd9, 12'sd1371}},
{{12'sd-2008, 12'sd1744, 13'sd-2070}, {12'sd1161, 13'sd-2581, 10'sd413}, {13'sd-2251, 12'sd-1374, 10'sd-289}},
{{12'sd-1747, 11'sd-703, 12'sd-1957}, {12'sd-1040, 13'sd2130, 11'sd-977}, {11'sd533, 12'sd-1466, 13'sd2181}},
{{13'sd-4069, 11'sd657, 6'sd18}, {13'sd-3448, 13'sd-2118, 13'sd3084}, {13'sd-3286, 12'sd-1636, 12'sd1074}},
{{12'sd-1191, 13'sd2632, 11'sd-980}, {13'sd-2384, 12'sd-1988, 13'sd2946}, {12'sd1440, 13'sd-3078, 9'sd143}},
{{9'sd223, 12'sd-1397, 12'sd1785}, {11'sd-675, 12'sd1799, 12'sd1063}, {13'sd2557, 13'sd2344, 12'sd-1106}},
{{13'sd-2261, 12'sd1061, 13'sd-2484}, {12'sd1220, 12'sd1543, 12'sd1979}, {11'sd-574, 4'sd5, 9'sd-145}},
{{12'sd1510, 13'sd-2544, 13'sd-2381}, {13'sd2586, 8'sd-114, 12'sd1331}, {12'sd1457, 10'sd320, 13'sd-2171}},
{{13'sd-2504, 12'sd1241, 9'sd246}, {11'sd927, 12'sd1772, 12'sd1596}, {13'sd3018, 11'sd893, 13'sd2592}},
{{11'sd799, 12'sd-1678, 11'sd-712}, {5'sd-8, 13'sd-2202, 13'sd2418}, {13'sd-2082, 9'sd-252, 13'sd2136}},
{{13'sd2361, 11'sd966, 13'sd-2476}, {13'sd-2145, 12'sd1349, 11'sd942}, {11'sd-531, 13'sd-2207, 9'sd163}},
{{13'sd-2126, 13'sd2608, 13'sd2751}, {13'sd2261, 12'sd1195, 12'sd1743}, {13'sd2112, 12'sd1358, 8'sd-104}},
{{13'sd-2681, 10'sd415, 13'sd2230}, {5'sd13, 12'sd1313, 13'sd2095}, {12'sd1231, 12'sd1108, 12'sd-1427}},
{{12'sd-1338, 11'sd-828, 13'sd2152}, {11'sd561, 11'sd-989, 11'sd-568}, {11'sd519, 12'sd-1269, 13'sd-2428}},
{{12'sd1203, 13'sd-2177, 12'sd1811}, {12'sd1348, 7'sd-47, 11'sd-816}, {11'sd-1014, 12'sd-1514, 13'sd2152}},
{{13'sd3092, 12'sd1696, 12'sd-1766}, {11'sd-517, 11'sd-647, 11'sd879}, {12'sd-1234, 13'sd-2218, 12'sd1553}},
{{7'sd45, 12'sd1935, 11'sd703}, {13'sd-3504, 13'sd-2500, 11'sd726}, {12'sd-1930, 12'sd1619, 11'sd-631}},
{{13'sd-2886, 11'sd-628, 11'sd887}, {13'sd-2271, 11'sd-649, 12'sd-1872}, {11'sd848, 10'sd-504, 13'sd2708}},
{{13'sd3670, 13'sd2203, 12'sd-1555}, {13'sd2080, 13'sd2908, 10'sd-442}, {10'sd326, 11'sd-866, 11'sd-527}},
{{13'sd-2473, 11'sd655, 11'sd808}, {11'sd622, 13'sd2607, 12'sd1197}, {12'sd-1085, 11'sd-748, 13'sd-2258}},
{{8'sd-125, 10'sd-466, 11'sd717}, {12'sd-1185, 13'sd2377, 12'sd1628}, {12'sd-1320, 13'sd2495, 11'sd-618}},
{{13'sd2413, 11'sd-936, 9'sd-244}, {12'sd1266, 12'sd1063, 13'sd2052}, {10'sd-352, 13'sd2552, 13'sd2438}},
{{11'sd928, 10'sd413, 13'sd2460}, {13'sd-2316, 7'sd-60, 13'sd-2060}, {11'sd-641, 13'sd-2333, 12'sd-1626}},
{{12'sd1544, 12'sd-1939, 13'sd2107}, {13'sd2658, 11'sd-930, 13'sd-2097}, {12'sd1077, 12'sd-1084, 8'sd73}},
{{8'sd-91, 12'sd1985, 13'sd-2647}, {12'sd1872, 11'sd-917, 13'sd-2528}, {11'sd591, 12'sd1892, 12'sd-1767}},
{{13'sd-2353, 13'sd-2629, 12'sd-1835}, {13'sd2361, 13'sd-2122, 12'sd1092}, {12'sd-2004, 12'sd2031, 11'sd-987}},
{{13'sd-2143, 12'sd1701, 12'sd1694}, {13'sd3110, 10'sd497, 11'sd847}, {7'sd53, 9'sd-180, 11'sd-864}},
{{13'sd2105, 11'sd-890, 12'sd-1601}, {13'sd2636, 12'sd-1324, 8'sd97}, {12'sd1863, 13'sd2322, 12'sd1754}},
{{12'sd1874, 12'sd-1637, 12'sd1418}, {8'sd105, 13'sd2550, 11'sd-757}, {11'sd-974, 12'sd-2015, 13'sd-2631}},
{{11'sd797, 11'sd991, 9'sd162}, {12'sd-1108, 13'sd2314, 13'sd-2137}, {13'sd-2213, 10'sd-488, 10'sd426}},
{{12'sd1258, 12'sd-1751, 12'sd1179}, {12'sd1442, 8'sd-74, 13'sd-2236}, {11'sd-807, 9'sd178, 13'sd-2865}},
{{9'sd-213, 10'sd305, 13'sd2290}, {11'sd822, 13'sd2401, 13'sd2671}, {12'sd-1739, 10'sd-453, 13'sd2601}},
{{12'sd-1285, 11'sd-629, 10'sd-437}, {12'sd-1752, 7'sd62, 7'sd-36}, {11'sd969, 11'sd627, 12'sd1830}},
{{8'sd94, 12'sd1101, 10'sd-340}, {12'sd-1253, 12'sd1332, 12'sd-1880}, {6'sd-27, 9'sd-163, 9'sd232}},
{{11'sd688, 12'sd-1497, 6'sd-30}, {10'sd313, 12'sd-1032, 9'sd-178}, {13'sd-3267, 13'sd2820, 13'sd2922}},
{{13'sd-2803, 12'sd-1978, 13'sd-2558}, {11'sd-516, 11'sd-718, 13'sd2258}, {12'sd2008, 8'sd104, 13'sd3117}},
{{13'sd2359, 13'sd2845, 10'sd345}, {10'sd293, 11'sd588, 12'sd-1622}, {13'sd2184, 11'sd-597, 9'sd137}},
{{13'sd-2655, 12'sd1103, 12'sd-1457}, {11'sd571, 6'sd31, 13'sd-2295}, {12'sd-2002, 11'sd-879, 12'sd-1521}},
{{12'sd1417, 11'sd-820, 10'sd-293}, {13'sd2866, 12'sd-1756, 13'sd-2102}, {10'sd278, 11'sd-892, 12'sd1716}},
{{12'sd1291, 12'sd-1644, 11'sd728}, {12'sd1072, 13'sd-2767, 13'sd-2905}, {11'sd-856, 11'sd-595, 9'sd-222}},
{{9'sd197, 12'sd-1865, 6'sd-18}, {10'sd504, 12'sd-1449, 11'sd-634}, {8'sd121, 13'sd2137, 12'sd-1429}},
{{10'sd443, 13'sd2574, 11'sd684}, {12'sd-1428, 11'sd948, 12'sd1492}, {9'sd-143, 12'sd1155, 12'sd1631}},
{{13'sd3153, 13'sd-2488, 13'sd2066}, {12'sd-1853, 13'sd-2638, 12'sd1248}, {13'sd3049, 13'sd-2078, 12'sd1121}},
{{10'sd-411, 13'sd-2221, 10'sd-377}, {12'sd1960, 12'sd-1110, 11'sd-524}, {13'sd-2301, 13'sd-2774, 12'sd1773}},
{{11'sd-868, 11'sd593, 11'sd-780}, {11'sd590, 12'sd1145, 12'sd1629}, {13'sd-3104, 12'sd1200, 12'sd-1761}},
{{12'sd-1434, 10'sd-477, 13'sd-2703}, {13'sd-2283, 13'sd-2202, 11'sd-894}, {12'sd1489, 12'sd1268, 12'sd1029}},
{{11'sd-807, 11'sd-865, 12'sd1807}, {11'sd-1016, 12'sd-1447, 12'sd1198}, {12'sd1904, 13'sd-2713, 13'sd-2304}},
{{13'sd3107, 12'sd-1375, 13'sd3029}, {11'sd-526, 12'sd-1750, 9'sd144}, {12'sd2006, 12'sd-1739, 9'sd-180}},
{{12'sd1036, 12'sd1417, 12'sd-1495}, {11'sd879, 10'sd439, 12'sd-1573}, {13'sd-2364, 12'sd1439, 12'sd-1758}},
{{13'sd-2980, 13'sd-2340, 10'sd-467}, {10'sd418, 11'sd-709, 9'sd-158}, {12'sd-1354, 12'sd-1334, 13'sd3067}}},
{
{{12'sd1172, 13'sd-3041, 12'sd-1559}, {13'sd-2368, 8'sd93, 13'sd-2268}, {13'sd-2835, 13'sd-2109, 11'sd669}},
{{13'sd3119, 12'sd1130, 12'sd1239}, {12'sd-1396, 13'sd-2131, 13'sd2183}, {12'sd-1364, 12'sd-1236, 13'sd2263}},
{{11'sd769, 12'sd1976, 9'sd-159}, {13'sd2220, 12'sd-1849, 11'sd795}, {10'sd390, 12'sd-1182, 13'sd-2806}},
{{13'sd-2538, 12'sd-1795, 9'sd-157}, {11'sd809, 13'sd-3106, 10'sd-452}, {13'sd-2844, 8'sd109, 11'sd-552}},
{{7'sd63, 11'sd783, 13'sd-2968}, {11'sd-523, 12'sd-1297, 9'sd-161}, {12'sd2008, 11'sd616, 7'sd51}},
{{10'sd266, 11'sd640, 13'sd-2760}, {11'sd-991, 13'sd-2295, 10'sd258}, {8'sd-92, 10'sd-443, 10'sd-295}},
{{12'sd1364, 12'sd1931, 11'sd-882}, {12'sd-1090, 12'sd-1731, 12'sd-1174}, {11'sd-696, 13'sd-3038, 9'sd-241}},
{{12'sd1832, 10'sd-473, 13'sd2671}, {11'sd-780, 13'sd-2590, 12'sd1308}, {13'sd-3001, 12'sd1065, 12'sd-1155}},
{{12'sd-1152, 12'sd-1599, 12'sd1591}, {13'sd-2577, 11'sd651, 10'sd-402}, {10'sd-436, 11'sd-859, 13'sd-2123}},
{{12'sd-2008, 11'sd977, 7'sd-34}, {12'sd1087, 12'sd-1437, 12'sd-1314}, {13'sd-2152, 12'sd1158, 9'sd130}},
{{13'sd2403, 11'sd-927, 13'sd2358}, {12'sd1192, 12'sd-1477, 13'sd2447}, {12'sd-1093, 12'sd1774, 12'sd1542}},
{{12'sd-1709, 12'sd1503, 11'sd-719}, {9'sd187, 9'sd141, 12'sd-1835}, {11'sd-767, 13'sd-2224, 13'sd2257}},
{{11'sd993, 11'sd-740, 12'sd1266}, {13'sd2504, 14'sd-4278, 13'sd-2317}, {12'sd-1807, 14'sd-5367, 14'sd-4670}},
{{10'sd321, 11'sd709, 12'sd-1819}, {10'sd-421, 12'sd-1278, 12'sd-1384}, {12'sd-1756, 11'sd-807, 10'sd-409}},
{{12'sd-1197, 9'sd-188, 12'sd-1119}, {10'sd-331, 11'sd-571, 12'sd-1837}, {12'sd-1687, 12'sd-1420, 12'sd1703}},
{{12'sd1399, 13'sd2372, 13'sd3150}, {9'sd149, 13'sd3105, 12'sd1135}, {12'sd1812, 12'sd-2031, 12'sd-1440}},
{{10'sd369, 12'sd-1268, 10'sd271}, {12'sd-1156, 12'sd1372, 13'sd-2441}, {11'sd-521, 10'sd314, 9'sd-202}},
{{13'sd-3670, 9'sd136, 13'sd2239}, {12'sd-1322, 12'sd-1389, 12'sd-1744}, {13'sd-2521, 10'sd-463, 11'sd-941}},
{{11'sd-591, 12'sd-1467, 12'sd1120}, {11'sd953, 8'sd-100, 12'sd1630}, {10'sd-287, 13'sd2348, 13'sd-2500}},
{{12'sd1830, 8'sd108, 12'sd1189}, {12'sd1990, 12'sd1807, 12'sd1593}, {12'sd1057, 12'sd1708, 11'sd941}},
{{12'sd1573, 12'sd1522, 12'sd1722}, {12'sd1552, 10'sd328, 12'sd1373}, {11'sd803, 13'sd2638, 12'sd1800}},
{{11'sd-912, 13'sd-2464, 12'sd-1413}, {13'sd-2217, 12'sd-1876, 12'sd-1415}, {11'sd-674, 13'sd-2809, 10'sd446}},
{{13'sd-2836, 13'sd-2230, 8'sd92}, {12'sd-1995, 11'sd821, 11'sd866}, {11'sd728, 12'sd-1979, 13'sd-2496}},
{{12'sd-1659, 10'sd-325, 12'sd-1376}, {8'sd-112, 12'sd1970, 12'sd1948}, {13'sd-2304, 13'sd2659, 12'sd-1560}},
{{13'sd-2305, 10'sd301, 9'sd222}, {13'sd-2261, 8'sd124, 12'sd-1824}, {11'sd-615, 11'sd-700, 13'sd3147}},
{{12'sd-1469, 8'sd65, 12'sd1388}, {11'sd920, 9'sd254, 12'sd-1574}, {11'sd-981, 11'sd873, 13'sd2286}},
{{13'sd-2496, 7'sd-55, 13'sd-2425}, {12'sd-1731, 10'sd368, 11'sd-1005}, {13'sd2228, 12'sd1844, 11'sd835}},
{{10'sd328, 12'sd1477, 11'sd698}, {11'sd1014, 9'sd-235, 12'sd-1059}, {11'sd735, 10'sd-435, 13'sd-2663}},
{{11'sd-989, 11'sd519, 9'sd-164}, {13'sd2591, 12'sd-1852, 11'sd974}, {12'sd1256, 9'sd-147, 13'sd2537}},
{{12'sd2021, 10'sd-316, 12'sd-1831}, {13'sd-2124, 12'sd-1999, 11'sd-878}, {13'sd-2222, 13'sd2733, 12'sd-1674}},
{{12'sd-1436, 13'sd2217, 13'sd2095}, {9'sd167, 13'sd3333, 13'sd2849}, {13'sd-2132, 13'sd2921, 11'sd-601}},
{{13'sd-2549, 11'sd758, 13'sd2319}, {11'sd940, 10'sd451, 13'sd2438}, {12'sd-1617, 12'sd1271, 13'sd2284}},
{{11'sd-766, 13'sd2117, 11'sd-514}, {12'sd-1813, 11'sd-831, 12'sd1491}, {12'sd1218, 12'sd1657, 11'sd736}},
{{11'sd-813, 10'sd-350, 7'sd43}, {11'sd732, 13'sd2051, 13'sd2640}, {12'sd-1559, 13'sd2550, 12'sd1352}},
{{12'sd1865, 13'sd2173, 11'sd542}, {13'sd-2331, 13'sd-2368, 11'sd-819}, {13'sd-2758, 11'sd571, 9'sd187}},
{{11'sd777, 13'sd2837, 12'sd1234}, {13'sd-2370, 13'sd2740, 12'sd-1459}, {13'sd2235, 12'sd-1347, 12'sd-1858}},
{{12'sd-1890, 12'sd1998, 12'sd1192}, {10'sd-475, 12'sd1387, 12'sd-1355}, {12'sd-1387, 12'sd-1344, 12'sd1663}},
{{13'sd2337, 12'sd-1353, 11'sd878}, {12'sd-1615, 12'sd2010, 11'sd711}, {13'sd2760, 13'sd-2397, 12'sd1833}},
{{9'sd222, 13'sd2505, 11'sd-914}, {12'sd-1233, 13'sd-2770, 13'sd-2742}, {13'sd-2537, 13'sd2535, 12'sd1747}},
{{11'sd944, 11'sd844, 13'sd2427}, {13'sd-2566, 13'sd2672, 13'sd-2430}, {12'sd-1664, 12'sd-1805, 8'sd93}},
{{9'sd-198, 11'sd-725, 13'sd-2905}, {11'sd519, 12'sd-1939, 12'sd-1058}, {12'sd2020, 11'sd-874, 11'sd705}},
{{13'sd2377, 12'sd1863, 13'sd2451}, {8'sd120, 12'sd1119, 12'sd2011}, {13'sd-2049, 11'sd-939, 13'sd-2070}},
{{11'sd908, 11'sd-952, 11'sd-637}, {9'sd130, 13'sd-2733, 11'sd697}, {12'sd1612, 12'sd1499, 10'sd-315}},
{{12'sd-1184, 10'sd446, 12'sd1886}, {13'sd-2380, 13'sd3025, 10'sd-450}, {12'sd-2043, 9'sd130, 9'sd131}},
{{12'sd-1288, 12'sd1357, 12'sd-1414}, {11'sd1018, 12'sd1946, 11'sd-853}, {9'sd183, 13'sd-2146, 12'sd-1437}},
{{12'sd-1147, 13'sd2432, 12'sd-1261}, {9'sd-255, 11'sd893, 12'sd1548}, {12'sd-1253, 11'sd-832, 12'sd1412}},
{{12'sd1947, 13'sd2559, 10'sd-309}, {11'sd765, 11'sd-780, 8'sd112}, {12'sd-1266, 13'sd2523, 13'sd2208}},
{{14'sd4432, 12'sd1355, 13'sd3044}, {11'sd-833, 12'sd-1558, 13'sd2542}, {11'sd-524, 11'sd512, 11'sd863}},
{{13'sd-2959, 12'sd1251, 8'sd-86}, {13'sd-4001, 13'sd2264, 11'sd850}, {12'sd-1653, 12'sd1408, 9'sd-157}},
{{11'sd-752, 12'sd1786, 12'sd-1113}, {13'sd-3706, 10'sd-433, 12'sd-1628}, {12'sd1594, 10'sd422, 10'sd426}},
{{12'sd1317, 12'sd1212, 12'sd-2036}, {12'sd2036, 12'sd1755, 12'sd-1956}, {13'sd2521, 12'sd-1480, 13'sd2158}},
{{11'sd926, 13'sd2131, 10'sd344}, {13'sd2075, 10'sd315, 11'sd-957}, {12'sd-1313, 7'sd34, 13'sd-2178}},
{{12'sd1720, 11'sd675, 12'sd-1978}, {12'sd-1094, 11'sd-866, 13'sd-2137}, {12'sd1364, 9'sd-235, 12'sd1606}},
{{11'sd-621, 11'sd-778, 12'sd1763}, {13'sd-3038, 11'sd-640, 13'sd2521}, {13'sd-2696, 10'sd259, 12'sd-1880}},
{{11'sd734, 11'sd-586, 11'sd-602}, {13'sd-2095, 10'sd431, 12'sd1081}, {13'sd-3760, 9'sd138, 13'sd-3855}},
{{11'sd-770, 11'sd1000, 11'sd-791}, {13'sd2456, 12'sd-1617, 12'sd-1581}, {13'sd2170, 8'sd-96, 12'sd1968}},
{{12'sd1543, 13'sd2136, 13'sd2118}, {8'sd-98, 12'sd1772, 11'sd-540}, {13'sd-2556, 12'sd1538, 11'sd533}},
{{13'sd3781, 11'sd858, 13'sd-2391}, {12'sd1565, 11'sd-846, 12'sd1179}, {12'sd-1247, 10'sd475, 13'sd-2462}},
{{13'sd2670, 12'sd-1630, 12'sd-1662}, {13'sd-2430, 12'sd-1601, 12'sd1888}, {6'sd-26, 12'sd-1629, 13'sd2463}},
{{13'sd3995, 11'sd798, 10'sd-361}, {12'sd1082, 13'sd-2128, 12'sd-1860}, {11'sd818, 9'sd182, 10'sd342}},
{{12'sd-1773, 10'sd413, 12'sd-1822}, {12'sd1928, 8'sd-126, 11'sd892}, {13'sd-2271, 13'sd2590, 13'sd2507}},
{{10'sd431, 11'sd995, 12'sd1885}, {13'sd-3054, 13'sd2282, 12'sd1988}, {11'sd-992, 12'sd-2028, 12'sd1443}},
{{12'sd1067, 13'sd2848, 11'sd567}, {12'sd-1092, 12'sd-1541, 10'sd-347}, {12'sd-1215, 12'sd1161, 7'sd39}},
{{13'sd2223, 11'sd-582, 9'sd-254}, {10'sd377, 10'sd-487, 10'sd272}, {6'sd-24, 13'sd-2241, 12'sd1513}}},
{
{{9'sd200, 12'sd-1725, 11'sd630}, {11'sd-743, 9'sd-146, 9'sd243}, {12'sd-1616, 8'sd75, 10'sd-302}},
{{12'sd-1990, 12'sd1041, 12'sd1301}, {12'sd1106, 11'sd794, 10'sd264}, {8'sd-126, 12'sd1523, 12'sd-1524}},
{{7'sd62, 13'sd-2999, 13'sd-3425}, {12'sd-1360, 12'sd-1091, 9'sd-144}, {13'sd2552, 9'sd-210, 10'sd492}},
{{9'sd184, 12'sd1136, 12'sd1853}, {13'sd2241, 10'sd267, 11'sd-638}, {13'sd2717, 13'sd3085, 13'sd2092}},
{{13'sd2421, 11'sd-598, 11'sd-552}, {13'sd-2517, 12'sd-1099, 10'sd-370}, {11'sd606, 10'sd-383, 12'sd1341}},
{{13'sd2199, 10'sd-289, 10'sd-335}, {12'sd-1783, 13'sd2115, 12'sd1282}, {12'sd1129, 12'sd-1712, 11'sd-746}},
{{12'sd-1880, 12'sd-1395, 10'sd-403}, {13'sd-2272, 10'sd-448, 12'sd-1501}, {13'sd-2074, 11'sd-938, 13'sd2421}},
{{12'sd1264, 12'sd-1434, 13'sd-2751}, {13'sd2129, 11'sd973, 13'sd2123}, {11'sd-534, 11'sd-654, 12'sd1796}},
{{8'sd89, 12'sd1136, 13'sd-2491}, {12'sd1963, 11'sd-712, 12'sd1890}, {11'sd-689, 12'sd-1978, 13'sd-3533}},
{{12'sd1052, 12'sd1248, 12'sd-1355}, {12'sd1488, 11'sd675, 13'sd-2314}, {13'sd-2578, 12'sd1289, 13'sd-2414}},
{{13'sd2287, 12'sd-1245, 12'sd-1603}, {13'sd2118, 12'sd-1905, 7'sd-50}, {11'sd-700, 11'sd851, 12'sd1671}},
{{11'sd-588, 12'sd1747, 13'sd-2253}, {9'sd-198, 12'sd1035, 11'sd-642}, {12'sd1078, 7'sd-59, 10'sd-485}},
{{13'sd-3267, 12'sd-1423, 9'sd150}, {13'sd-2722, 10'sd330, 12'sd-1234}, {10'sd460, 12'sd1101, 13'sd-2236}},
{{8'sd-109, 13'sd-2731, 12'sd-1899}, {9'sd-149, 10'sd-337, 12'sd1854}, {12'sd1711, 13'sd-2579, 11'sd-1021}},
{{12'sd1611, 13'sd2114, 11'sd954}, {13'sd-3245, 10'sd-309, 13'sd-2577}, {12'sd1792, 12'sd-1815, 11'sd937}},
{{9'sd203, 12'sd1412, 13'sd2283}, {12'sd1861, 10'sd339, 13'sd-2136}, {12'sd-1430, 13'sd-2088, 12'sd-2019}},
{{7'sd40, 13'sd2116, 12'sd1937}, {13'sd2472, 11'sd625, 11'sd666}, {10'sd-402, 11'sd750, 10'sd-364}},
{{12'sd1222, 11'sd657, 10'sd425}, {11'sd539, 12'sd1076, 13'sd-2490}, {13'sd2285, 11'sd837, 13'sd-3328}},
{{9'sd-207, 12'sd-1592, 8'sd107}, {11'sd712, 10'sd-356, 12'sd-1945}, {12'sd-1602, 11'sd809, 9'sd220}},
{{10'sd-384, 13'sd2257, 13'sd2314}, {11'sd979, 11'sd-609, 11'sd936}, {12'sd1271, 13'sd-2657, 12'sd1314}},
{{13'sd-2532, 13'sd-2297, 12'sd1404}, {11'sd783, 12'sd1801, 12'sd-1271}, {8'sd-64, 9'sd196, 10'sd-346}},
{{12'sd1439, 11'sd580, 10'sd451}, {11'sd889, 11'sd565, 8'sd-81}, {12'sd1566, 12'sd1062, 12'sd1700}},
{{12'sd-1350, 12'sd-1500, 13'sd-2351}, {11'sd642, 12'sd-1657, 11'sd-811}, {11'sd892, 6'sd-19, 13'sd-2736}},
{{13'sd2136, 12'sd-1690, 8'sd113}, {13'sd-2307, 11'sd953, 12'sd-1046}, {13'sd2151, 12'sd1443, 11'sd611}},
{{8'sd-110, 12'sd-1983, 12'sd1055}, {10'sd-343, 12'sd-1191, 12'sd-1360}, {12'sd-1164, 12'sd-1958, 12'sd1033}},
{{12'sd1716, 11'sd576, 11'sd665}, {13'sd-2536, 13'sd2287, 12'sd1881}, {9'sd187, 12'sd1393, 12'sd-1458}},
{{12'sd-1165, 12'sd1820, 12'sd1942}, {11'sd-640, 11'sd-728, 13'sd2058}, {13'sd2694, 13'sd2740, 13'sd-2352}},
{{12'sd1278, 10'sd349, 9'sd136}, {11'sd592, 12'sd1778, 12'sd1694}, {12'sd-1625, 12'sd-1780, 13'sd2965}},
{{12'sd1753, 13'sd-2912, 11'sd591}, {11'sd-630, 10'sd-429, 12'sd-1948}, {11'sd957, 13'sd-2364, 10'sd484}},
{{13'sd2870, 10'sd-501, 12'sd-1576}, {13'sd-2547, 13'sd-2666, 12'sd1134}, {12'sd1332, 12'sd1423, 9'sd131}},
{{12'sd1723, 11'sd595, 13'sd2416}, {13'sd3702, 12'sd1599, 13'sd-3959}, {10'sd401, 13'sd2447, 12'sd-1573}},
{{12'sd-1523, 9'sd-192, 10'sd-361}, {12'sd1081, 13'sd2101, 13'sd2147}, {13'sd2193, 13'sd-2520, 4'sd-6}},
{{11'sd830, 11'sd-891, 3'sd-2}, {12'sd1571, 12'sd-1032, 13'sd-2365}, {10'sd-266, 13'sd2293, 11'sd616}},
{{13'sd-2978, 13'sd-2701, 11'sd-845}, {11'sd964, 10'sd-449, 12'sd-1093}, {10'sd-330, 12'sd1069, 12'sd1285}},
{{10'sd438, 12'sd-1507, 11'sd893}, {12'sd1602, 13'sd-2081, 11'sd-668}, {12'sd1257, 13'sd2080, 13'sd2368}},
{{11'sd-891, 12'sd-1150, 11'sd-753}, {11'sd832, 11'sd768, 11'sd-692}, {13'sd-2359, 12'sd1862, 12'sd1069}},
{{10'sd-473, 12'sd1425, 13'sd2625}, {13'sd-2095, 13'sd2338, 13'sd2460}, {12'sd-2025, 9'sd-225, 8'sd84}},
{{9'sd-207, 12'sd1978, 12'sd-1680}, {11'sd-926, 12'sd-1596, 11'sd-982}, {12'sd-1347, 13'sd2605, 9'sd-255}},
{{13'sd-2160, 11'sd-748, 12'sd1388}, {12'sd1071, 13'sd-2955, 11'sd788}, {11'sd838, 11'sd573, 11'sd844}},
{{13'sd-2380, 10'sd327, 13'sd-2691}, {12'sd-1449, 10'sd-314, 12'sd-1312}, {13'sd2511, 10'sd-315, 13'sd2517}},
{{13'sd-3282, 5'sd-13, 12'sd-1316}, {12'sd1749, 13'sd-2642, 13'sd2119}, {13'sd-3851, 11'sd-606, 10'sd357}},
{{12'sd-1322, 12'sd1199, 11'sd973}, {11'sd900, 12'sd-1229, 13'sd-2877}, {13'sd-2809, 13'sd-3638, 13'sd-2965}},
{{13'sd-3158, 12'sd-1604, 9'sd-144}, {13'sd-2833, 12'sd-1451, 13'sd3054}, {10'sd272, 13'sd-2185, 13'sd2267}},
{{9'sd-240, 10'sd-406, 11'sd-774}, {12'sd-1262, 11'sd573, 13'sd-2259}, {12'sd-1654, 11'sd-742, 10'sd-324}},
{{12'sd-1486, 12'sd-1037, 12'sd-1868}, {12'sd-1858, 12'sd-1036, 12'sd1278}, {13'sd-3035, 10'sd264, 12'sd-1777}},
{{12'sd1223, 12'sd1144, 12'sd-1647}, {12'sd1459, 13'sd2514, 13'sd-2461}, {12'sd1779, 11'sd-931, 9'sd-148}},
{{7'sd-55, 11'sd-1020, 9'sd-154}, {8'sd-108, 13'sd-2572, 12'sd-1289}, {11'sd-824, 12'sd1911, 12'sd-2019}},
{{13'sd-2697, 9'sd165, 13'sd-2761}, {12'sd-1325, 12'sd-1373, 13'sd2221}, {13'sd-2687, 13'sd-2577, 13'sd-3286}},
{{10'sd404, 13'sd2185, 13'sd2365}, {12'sd1406, 12'sd1300, 11'sd-577}, {13'sd3711, 6'sd-23, 13'sd2710}},
{{12'sd-1730, 8'sd80, 11'sd879}, {13'sd-2410, 8'sd-65, 13'sd-2331}, {13'sd2966, 12'sd-1097, 9'sd-151}},
{{11'sd831, 9'sd-211, 13'sd2171}, {4'sd5, 9'sd193, 11'sd-964}, {10'sd-477, 10'sd-497, 12'sd-1705}},
{{13'sd-2462, 13'sd-2455, 12'sd1407}, {12'sd-1509, 12'sd-1871, 12'sd1861}, {11'sd-745, 12'sd1257, 12'sd1965}},
{{12'sd-1379, 13'sd-2333, 12'sd1166}, {13'sd-2049, 10'sd-506, 12'sd1223}, {13'sd2969, 13'sd2393, 10'sd403}},
{{12'sd1819, 9'sd210, 12'sd1284}, {12'sd1309, 12'sd1636, 11'sd-938}, {12'sd-1611, 13'sd2151, 12'sd-1558}},
{{11'sd-529, 12'sd-1847, 12'sd1726}, {13'sd3156, 9'sd146, 10'sd400}, {7'sd-33, 10'sd-493, 12'sd1041}},
{{12'sd-1966, 11'sd890, 11'sd-623}, {11'sd894, 6'sd20, 13'sd2322}, {10'sd-373, 11'sd-677, 13'sd-2306}},
{{13'sd-2118, 13'sd-2942, 12'sd-1193}, {13'sd-2263, 7'sd-35, 12'sd-1088}, {11'sd-589, 12'sd1601, 13'sd2218}},
{{13'sd-2978, 13'sd2159, 13'sd-2133}, {11'sd604, 13'sd2597, 11'sd923}, {13'sd-2079, 11'sd601, 13'sd-2382}},
{{13'sd2545, 12'sd-1214, 12'sd-1400}, {12'sd1897, 12'sd-1201, 13'sd-2067}, {12'sd2002, 13'sd2134, 12'sd-1300}},
{{12'sd-1203, 13'sd-2311, 12'sd-1724}, {12'sd1191, 9'sd138, 13'sd-2579}, {13'sd2057, 12'sd-1914, 13'sd-3043}},
{{12'sd-1266, 13'sd-2240, 10'sd353}, {13'sd2526, 12'sd1445, 13'sd-2067}, {11'sd-993, 10'sd-445, 10'sd-409}},
{{11'sd-907, 12'sd1358, 12'sd-1103}, {10'sd347, 12'sd1647, 13'sd-2803}, {10'sd-444, 13'sd-2050, 7'sd-61}},
{{11'sd550, 11'sd-947, 13'sd-2510}, {12'sd1264, 10'sd368, 12'sd1364}, {12'sd1897, 12'sd1575, 12'sd-1040}},
{{13'sd-2395, 10'sd416, 12'sd-1730}, {10'sd-285, 12'sd-1788, 12'sd-2028}, {12'sd-1809, 12'sd1713, 13'sd-3006}}},
{
{{13'sd2479, 13'sd2128, 12'sd1384}, {12'sd-1394, 11'sd-867, 10'sd452}, {11'sd-896, 11'sd-866, 12'sd2034}},
{{11'sd-869, 13'sd2820, 3'sd3}, {10'sd-298, 12'sd-1353, 13'sd-2425}, {12'sd1944, 11'sd-836, 13'sd-2442}},
{{9'sd232, 10'sd-363, 10'sd-438}, {12'sd-1580, 13'sd2197, 9'sd-207}, {14'sd4152, 14'sd4191, 11'sd-772}},
{{11'sd-866, 10'sd349, 11'sd969}, {12'sd1960, 12'sd-1501, 12'sd-1244}, {13'sd2270, 12'sd1349, 10'sd-368}},
{{12'sd-1501, 13'sd2992, 13'sd2217}, {12'sd-1443, 13'sd-2475, 13'sd2928}, {11'sd781, 12'sd1854, 10'sd-326}},
{{13'sd2079, 9'sd224, 12'sd-1102}, {12'sd-1314, 11'sd-1018, 9'sd-226}, {13'sd2368, 12'sd1028, 13'sd-2419}},
{{13'sd2461, 11'sd-679, 13'sd2573}, {13'sd-2215, 11'sd-997, 12'sd-1345}, {12'sd-1397, 13'sd-3035, 10'sd372}},
{{12'sd1909, 10'sd-291, 13'sd3340}, {11'sd687, 13'sd-3128, 12'sd-1871}, {13'sd3081, 7'sd63, 8'sd95}},
{{12'sd1517, 13'sd-2455, 10'sd-467}, {13'sd3127, 12'sd-1948, 13'sd2600}, {10'sd-410, 13'sd2650, 11'sd592}},
{{11'sd652, 10'sd-474, 11'sd-880}, {9'sd-176, 12'sd-1936, 13'sd2680}, {12'sd1694, 8'sd-126, 9'sd-243}},
{{12'sd1358, 7'sd35, 12'sd-1237}, {13'sd2649, 11'sd-1003, 11'sd662}, {13'sd2270, 12'sd2014, 9'sd183}},
{{12'sd-1775, 13'sd2471, 7'sd34}, {10'sd294, 12'sd-1771, 12'sd-1538}, {12'sd-2023, 11'sd890, 12'sd-1045}},
{{13'sd-2062, 12'sd1648, 12'sd1106}, {13'sd-3751, 11'sd770, 13'sd-2633}, {12'sd-1980, 12'sd1926, 11'sd1016}},
{{13'sd2180, 11'sd-606, 12'sd-1431}, {12'sd1329, 11'sd-939, 13'sd2083}, {10'sd375, 10'sd-495, 11'sd915}},
{{11'sd-650, 13'sd-2519, 12'sd1109}, {13'sd2872, 12'sd-1101, 13'sd3247}, {9'sd158, 13'sd-2246, 13'sd3492}},
{{13'sd-2306, 7'sd-37, 12'sd-1801}, {12'sd-1184, 12'sd-1523, 13'sd-2416}, {11'sd769, 12'sd-1142, 11'sd-803}},
{{11'sd739, 12'sd-1129, 12'sd-1424}, {9'sd188, 13'sd-2135, 10'sd-373}, {12'sd-1504, 8'sd-104, 12'sd1840}},
{{11'sd597, 13'sd3992, 13'sd2999}, {13'sd2651, 12'sd1706, 14'sd4457}, {12'sd-1491, 12'sd1949, 13'sd3934}},
{{11'sd-968, 11'sd-581, 13'sd3022}, {13'sd3180, 12'sd-1491, 11'sd853}, {13'sd-2144, 12'sd1740, 12'sd-1839}},
{{7'sd54, 12'sd2038, 11'sd950}, {8'sd-88, 12'sd-1915, 11'sd-698}, {11'sd-540, 12'sd1186, 6'sd21}},
{{13'sd-3181, 8'sd-106, 9'sd-152}, {11'sd-556, 12'sd-2008, 12'sd1104}, {10'sd461, 12'sd1305, 10'sd-412}},
{{12'sd-1655, 13'sd-2440, 11'sd-752}, {13'sd2795, 12'sd-1937, 10'sd431}, {10'sd-477, 13'sd-2789, 11'sd809}},
{{12'sd-1665, 11'sd-911, 13'sd3113}, {9'sd-213, 10'sd-472, 12'sd-1215}, {13'sd2169, 10'sd-328, 12'sd-1186}},
{{11'sd800, 12'sd1705, 13'sd2353}, {13'sd2244, 13'sd-2151, 12'sd-1620}, {12'sd1778, 12'sd-1267, 12'sd-1254}},
{{12'sd1099, 12'sd-1935, 13'sd2306}, {13'sd2541, 12'sd-1843, 12'sd-1631}, {12'sd1251, 9'sd-247, 11'sd616}},
{{11'sd-961, 12'sd-1445, 12'sd1921}, {13'sd2237, 12'sd1165, 13'sd-2317}, {12'sd-1870, 12'sd1668, 12'sd1669}},
{{13'sd2517, 12'sd2018, 12'sd-2016}, {13'sd-2778, 11'sd806, 13'sd-2797}, {12'sd1953, 12'sd1123, 12'sd-1713}},
{{13'sd2341, 13'sd3605, 12'sd1910}, {11'sd-1010, 12'sd-1323, 12'sd-1261}, {13'sd-2571, 12'sd-1036, 10'sd428}},
{{13'sd-2352, 12'sd-1669, 12'sd1601}, {10'sd376, 13'sd-2535, 11'sd802}, {13'sd2174, 13'sd-2849, 11'sd-623}},
{{9'sd231, 13'sd-2382, 11'sd-625}, {8'sd-79, 8'sd-78, 12'sd-1452}, {13'sd-3271, 12'sd1121, 12'sd-2037}},
{{12'sd1198, 10'sd-399, 11'sd-946}, {13'sd-2491, 11'sd803, 11'sd735}, {13'sd-3603, 11'sd-726, 12'sd-1179}},
{{12'sd-1331, 10'sd-362, 13'sd2880}, {13'sd2826, 13'sd2654, 8'sd-88}, {12'sd1029, 12'sd1636, 13'sd2811}},
{{12'sd-1270, 13'sd2768, 9'sd-136}, {9'sd183, 13'sd-2396, 11'sd727}, {11'sd-699, 12'sd1363, 10'sd504}},
{{3'sd-2, 9'sd-223, 11'sd-766}, {13'sd-2240, 12'sd1043, 11'sd620}, {12'sd1402, 12'sd1517, 13'sd-2069}},
{{12'sd1751, 8'sd124, 12'sd1286}, {11'sd740, 13'sd-2998, 11'sd-551}, {13'sd-2163, 12'sd-1865, 13'sd-2196}},
{{10'sd-486, 12'sd-1042, 10'sd304}, {12'sd-1910, 11'sd589, 12'sd1658}, {12'sd-1696, 11'sd-843, 12'sd1806}},
{{8'sd94, 12'sd1450, 13'sd2183}, {13'sd-2403, 13'sd-3228, 12'sd1604}, {7'sd-53, 13'sd-2130, 13'sd-2428}},
{{12'sd1519, 13'sd-2109, 10'sd472}, {11'sd672, 9'sd245, 12'sd-1471}, {11'sd606, 11'sd603, 12'sd-1381}},
{{12'sd-1940, 12'sd1422, 13'sd2081}, {13'sd-2952, 12'sd-1177, 11'sd-1003}, {12'sd-1227, 11'sd644, 13'sd-2228}},
{{11'sd-622, 13'sd-2337, 12'sd-1231}, {11'sd742, 11'sd965, 12'sd1076}, {13'sd-2578, 10'sd361, 12'sd-1195}},
{{13'sd2326, 12'sd-1594, 11'sd838}, {13'sd3593, 12'sd-1775, 12'sd1222}, {12'sd1560, 9'sd134, 9'sd178}},
{{11'sd-520, 12'sd1361, 12'sd1590}, {13'sd-2450, 12'sd-1571, 12'sd-1219}, {12'sd1467, 11'sd-578, 11'sd532}},
{{7'sd60, 12'sd1045, 12'sd1456}, {12'sd-1558, 12'sd1869, 12'sd1076}, {13'sd2733, 9'sd-177, 11'sd-933}},
{{11'sd807, 13'sd-2296, 9'sd-171}, {13'sd-2060, 9'sd-130, 12'sd1571}, {12'sd-1564, 11'sd-522, 11'sd846}},
{{13'sd-2229, 11'sd706, 12'sd-1164}, {8'sd120, 13'sd-3349, 12'sd1437}, {9'sd-182, 10'sd308, 10'sd-450}},
{{12'sd1870, 13'sd2760, 12'sd-1954}, {11'sd612, 11'sd-569, 11'sd679}, {13'sd2572, 12'sd1846, 13'sd-2603}},
{{12'sd2010, 11'sd-817, 11'sd-528}, {13'sd-2049, 7'sd54, 11'sd-519}, {9'sd-243, 13'sd2366, 11'sd1023}},
{{8'sd-71, 11'sd551, 10'sd-315}, {12'sd1729, 12'sd-2023, 12'sd1860}, {12'sd-1244, 9'sd-218, 12'sd-1495}},
{{12'sd-1517, 12'sd-1120, 11'sd-560}, {13'sd2064, 13'sd-2670, 11'sd921}, {12'sd1217, 13'sd2474, 10'sd338}},
{{12'sd1760, 12'sd-1260, 12'sd1893}, {13'sd2405, 10'sd504, 12'sd1467}, {13'sd3274, 13'sd2343, 14'sd5204}},
{{12'sd-1344, 5'sd14, 13'sd2135}, {12'sd1175, 11'sd-858, 12'sd1959}, {11'sd572, 12'sd1694, 12'sd1170}},
{{11'sd-706, 11'sd872, 13'sd2746}, {11'sd-635, 12'sd1129, 11'sd713}, {12'sd1067, 13'sd-2331, 13'sd-2904}},
{{12'sd-1037, 11'sd729, 9'sd216}, {13'sd-3010, 12'sd-1465, 13'sd-2237}, {13'sd-3327, 13'sd-2062, 12'sd1348}},
{{10'sd-270, 7'sd-33, 12'sd2022}, {12'sd-1294, 11'sd-884, 12'sd-1857}, {11'sd554, 12'sd-1509, 12'sd1072}},
{{10'sd497, 12'sd1253, 13'sd-3005}, {13'sd-2272, 11'sd-757, 10'sd-473}, {11'sd512, 12'sd-1372, 11'sd-876}},
{{11'sd742, 10'sd-358, 13'sd-2709}, {13'sd2085, 11'sd-885, 12'sd-1563}, {9'sd237, 11'sd591, 13'sd2493}},
{{11'sd693, 12'sd-1575, 13'sd2513}, {13'sd2621, 13'sd-2824, 10'sd-359}, {10'sd274, 8'sd85, 13'sd-2543}},
{{13'sd2049, 11'sd894, 12'sd-1986}, {13'sd3297, 11'sd806, 11'sd845}, {10'sd-290, 9'sd168, 11'sd567}},
{{10'sd-502, 12'sd1497, 12'sd-1716}, {13'sd-2572, 13'sd-3082, 12'sd-1601}, {11'sd-756, 12'sd-1704, 11'sd-941}},
{{7'sd-62, 11'sd971, 9'sd-250}, {11'sd810, 12'sd-1193, 12'sd-1910}, {13'sd-3812, 13'sd2310, 13'sd-2614}},
{{12'sd2018, 7'sd-48, 9'sd255}, {12'sd-1747, 13'sd2583, 9'sd-135}, {12'sd1793, 11'sd525, 12'sd1946}},
{{12'sd1841, 11'sd-948, 12'sd1855}, {13'sd-2101, 13'sd2094, 11'sd-882}, {12'sd1914, 12'sd-1736, 10'sd480}},
{{11'sd-684, 12'sd-1279, 11'sd698}, {12'sd-2011, 12'sd-1507, 12'sd-1102}, {11'sd-701, 13'sd-2481, 10'sd275}},
{{12'sd1933, 12'sd-1788, 11'sd819}, {13'sd-2165, 12'sd1175, 10'sd419}, {12'sd-1794, 13'sd2678, 11'sd-738}}},
{
{{13'sd2277, 5'sd15, 13'sd2328}, {13'sd-2104, 12'sd-1828, 11'sd-515}, {11'sd-1014, 10'sd411, 6'sd27}},
{{12'sd1339, 9'sd-191, 11'sd857}, {12'sd1328, 12'sd2003, 9'sd171}, {8'sd-101, 6'sd17, 9'sd-243}},
{{12'sd1246, 13'sd-2595, 12'sd1112}, {13'sd2089, 10'sd414, 13'sd2460}, {11'sd-971, 13'sd2214, 11'sd-901}},
{{12'sd1397, 13'sd2196, 12'sd1097}, {12'sd-1101, 12'sd-1825, 13'sd-2357}, {13'sd3219, 12'sd-1132, 13'sd2344}},
{{8'sd-104, 12'sd-1879, 11'sd-899}, {13'sd-2066, 13'sd2219, 10'sd377}, {12'sd-1452, 12'sd1407, 11'sd-943}},
{{12'sd-1629, 8'sd109, 12'sd-1395}, {13'sd-2150, 12'sd2039, 13'sd-2499}, {11'sd-689, 11'sd-704, 6'sd-31}},
{{11'sd-584, 11'sd1009, 12'sd-1117}, {12'sd-1807, 12'sd-1726, 10'sd-286}, {13'sd-3274, 13'sd-2564, 13'sd-2051}},
{{12'sd1837, 12'sd1711, 13'sd2529}, {12'sd2019, 11'sd652, 11'sd-814}, {10'sd397, 12'sd-1475, 13'sd-2186}},
{{11'sd877, 12'sd-1185, 13'sd2288}, {12'sd-2028, 13'sd2798, 8'sd-78}, {11'sd-933, 12'sd1390, 11'sd788}},
{{13'sd-2364, 13'sd2320, 13'sd2379}, {6'sd-25, 11'sd-995, 11'sd-757}, {12'sd-1792, 11'sd-576, 12'sd2047}},
{{12'sd1075, 13'sd2247, 12'sd-1395}, {12'sd1824, 11'sd-730, 10'sd365}, {11'sd-928, 12'sd-1142, 12'sd-1164}},
{{12'sd-1975, 5'sd10, 12'sd-1283}, {13'sd-2435, 12'sd-1135, 12'sd-1919}, {13'sd-2838, 11'sd-695, 12'sd1597}},
{{13'sd2285, 11'sd938, 13'sd3527}, {13'sd2942, 12'sd-1140, 13'sd2759}, {11'sd-512, 11'sd865, 13'sd-2429}},
{{11'sd-748, 12'sd2044, 10'sd-440}, {13'sd3016, 11'sd-876, 11'sd-562}, {13'sd-2742, 12'sd-1471, 13'sd2213}},
{{10'sd-275, 11'sd-549, 12'sd1195}, {12'sd1308, 13'sd-2519, 13'sd-2376}, {8'sd-100, 12'sd1994, 13'sd2683}},
{{13'sd-2461, 13'sd-2527, 10'sd385}, {11'sd-690, 13'sd-2642, 12'sd-1072}, {10'sd368, 12'sd1357, 13'sd2371}},
{{11'sd-791, 11'sd-868, 13'sd2452}, {9'sd159, 13'sd-2134, 13'sd-2098}, {13'sd-2578, 10'sd438, 13'sd-2069}},
{{11'sd-870, 10'sd495, 11'sd-762}, {12'sd-1677, 12'sd-1498, 6'sd23}, {12'sd-1476, 8'sd-109, 12'sd1957}},
{{13'sd2966, 12'sd1139, 12'sd-1608}, {9'sd162, 12'sd1308, 12'sd-1492}, {10'sd258, 13'sd-2311, 13'sd-2620}},
{{12'sd1871, 11'sd-765, 12'sd2019}, {12'sd1898, 10'sd-493, 12'sd-1834}, {11'sd-597, 13'sd-2493, 11'sd-884}},
{{13'sd-2759, 13'sd2171, 11'sd-922}, {12'sd-1519, 8'sd92, 10'sd-382}, {11'sd-733, 11'sd-770, 8'sd73}},
{{12'sd1984, 12'sd1177, 12'sd-1512}, {13'sd-2144, 10'sd489, 11'sd-685}, {12'sd-1856, 13'sd-2436, 12'sd1895}},
{{12'sd-1115, 12'sd1134, 11'sd684}, {12'sd-1335, 12'sd-1899, 6'sd23}, {11'sd-849, 12'sd-1416, 13'sd2523}},
{{13'sd-2975, 12'sd-1316, 12'sd1405}, {11'sd-603, 12'sd-1098, 11'sd694}, {12'sd1156, 11'sd-970, 12'sd1985}},
{{9'sd-197, 11'sd743, 12'sd-1240}, {11'sd541, 9'sd199, 13'sd2246}, {13'sd-2254, 11'sd835, 9'sd218}},
{{13'sd2090, 13'sd2499, 8'sd-104}, {12'sd-1432, 9'sd137, 12'sd-1471}, {13'sd-2330, 12'sd-1053, 13'sd2422}},
{{10'sd384, 11'sd520, 10'sd509}, {13'sd-2650, 13'sd-2335, 12'sd1690}, {10'sd-315, 12'sd-1198, 12'sd-1756}},
{{12'sd-1063, 13'sd2435, 12'sd1029}, {9'sd-128, 12'sd1847, 13'sd2091}, {12'sd1831, 12'sd-1734, 12'sd1429}},
{{12'sd-1849, 11'sd-876, 12'sd-1597}, {13'sd3041, 9'sd-139, 12'sd-1920}, {10'sd432, 13'sd-2141, 12'sd-1802}},
{{13'sd2637, 10'sd367, 13'sd-2395}, {12'sd1582, 13'sd-2423, 12'sd-1358}, {12'sd-1850, 13'sd2170, 13'sd2128}},
{{13'sd-3200, 12'sd-1315, 12'sd-1705}, {11'sd712, 13'sd-3917, 13'sd-3028}, {12'sd-1174, 10'sd-285, 11'sd-721}},
{{8'sd111, 13'sd-2400, 12'sd-1770}, {12'sd1890, 10'sd316, 12'sd1830}, {12'sd1058, 12'sd-1303, 10'sd287}},
{{12'sd1968, 12'sd-1790, 13'sd-2664}, {12'sd-1479, 13'sd2667, 12'sd1261}, {12'sd1266, 11'sd768, 11'sd657}},
{{12'sd1658, 11'sd893, 13'sd3335}, {12'sd1933, 12'sd1442, 12'sd-1105}, {12'sd-1475, 12'sd-1562, 12'sd1195}},
{{12'sd1687, 11'sd-925, 12'sd1392}, {12'sd-1716, 12'sd1276, 12'sd1612}, {12'sd-1040, 12'sd1839, 12'sd1754}},
{{12'sd-1475, 11'sd-515, 10'sd466}, {12'sd-1391, 11'sd737, 12'sd1697}, {11'sd939, 11'sd909, 13'sd-2080}},
{{11'sd830, 10'sd-469, 10'sd357}, {12'sd1621, 12'sd-1059, 13'sd-2129}, {12'sd1089, 2'sd-1, 12'sd-1616}},
{{12'sd1977, 13'sd2141, 13'sd2655}, {12'sd-1331, 13'sd-2511, 12'sd-1600}, {13'sd-2909, 6'sd-23, 13'sd-2489}},
{{13'sd2153, 13'sd2078, 13'sd2671}, {12'sd1771, 10'sd-302, 12'sd1469}, {13'sd2068, 12'sd-1105, 13'sd2195}},
{{10'sd509, 10'sd443, 12'sd1435}, {12'sd-1376, 8'sd-95, 10'sd-384}, {13'sd2153, 11'sd681, 12'sd1390}},
{{8'sd-119, 13'sd-2168, 13'sd2559}, {11'sd853, 8'sd-89, 13'sd3046}, {10'sd364, 12'sd-1902, 9'sd153}},
{{13'sd2500, 12'sd1469, 12'sd-1734}, {11'sd1010, 9'sd-156, 11'sd719}, {13'sd2738, 9'sd140, 12'sd-1485}},
{{12'sd-2012, 12'sd1982, 12'sd1707}, {12'sd1364, 12'sd-2012, 12'sd1844}, {12'sd1378, 5'sd13, 12'sd-2014}},
{{9'sd-169, 12'sd-1054, 12'sd1748}, {12'sd2031, 11'sd919, 13'sd-2598}, {11'sd-806, 11'sd-644, 12'sd-1054}},
{{13'sd-2156, 12'sd-1234, 13'sd2373}, {8'sd-72, 11'sd580, 8'sd111}, {11'sd-832, 10'sd333, 11'sd948}},
{{13'sd2081, 13'sd2798, 12'sd-1978}, {12'sd-1790, 10'sd477, 13'sd2536}, {7'sd-37, 10'sd-478, 12'sd-1437}},
{{12'sd-1510, 13'sd2330, 12'sd1555}, {12'sd-1192, 10'sd283, 12'sd1683}, {13'sd2185, 13'sd2101, 13'sd2616}},
{{10'sd-389, 10'sd498, 12'sd1962}, {11'sd-722, 13'sd2618, 13'sd-2556}, {13'sd-3149, 10'sd409, 10'sd374}},
{{12'sd1491, 12'sd1250, 11'sd-970}, {13'sd-2893, 10'sd267, 10'sd330}, {11'sd-644, 12'sd1346, 11'sd746}},
{{11'sd-774, 12'sd-1670, 11'sd680}, {13'sd-3415, 12'sd-1120, 13'sd-3091}, {13'sd-3329, 11'sd538, 13'sd-3277}},
{{12'sd1557, 12'sd1964, 11'sd526}, {10'sd-399, 13'sd-2274, 11'sd758}, {13'sd2594, 11'sd956, 11'sd-1009}},
{{13'sd2678, 12'sd1610, 11'sd932}, {11'sd976, 12'sd-1398, 11'sd674}, {13'sd2750, 12'sd-1534, 13'sd2861}},
{{13'sd2835, 13'sd-2075, 12'sd1142}, {10'sd-416, 11'sd576, 9'sd-198}, {12'sd-1654, 13'sd-2130, 12'sd1780}},
{{11'sd-823, 11'sd-719, 13'sd2552}, {10'sd-438, 9'sd173, 10'sd383}, {11'sd-761, 12'sd-1692, 9'sd-154}},
{{11'sd-669, 12'sd1124, 13'sd2523}, {12'sd1988, 13'sd-2682, 12'sd1208}, {13'sd2332, 13'sd2194, 12'sd1291}},
{{11'sd-845, 13'sd-2585, 13'sd2374}, {12'sd-1785, 12'sd-1104, 12'sd-2023}, {12'sd-1094, 11'sd-657, 12'sd-1178}},
{{12'sd1771, 11'sd-518, 11'sd-845}, {13'sd-2120, 12'sd-1610, 12'sd-1791}, {9'sd-185, 13'sd2209, 10'sd469}},
{{11'sd575, 10'sd431, 12'sd-1841}, {13'sd2533, 9'sd210, 12'sd-2031}, {12'sd-1661, 13'sd2681, 11'sd-996}},
{{12'sd1176, 12'sd1357, 12'sd-1616}, {10'sd455, 9'sd175, 12'sd1714}, {12'sd1405, 12'sd-1854, 8'sd-69}},
{{11'sd-550, 12'sd-1445, 13'sd2085}, {12'sd1189, 12'sd-1393, 12'sd1027}, {11'sd-769, 12'sd1597, 12'sd-1915}},
{{10'sd332, 7'sd63, 10'sd-405}, {12'sd-1805, 13'sd-2552, 12'sd1375}, {13'sd2311, 12'sd1723, 13'sd-2101}},
{{11'sd974, 10'sd289, 12'sd-1936}, {12'sd1619, 12'sd-1761, 13'sd-2574}, {8'sd-64, 13'sd-3329, 13'sd-2209}},
{{10'sd-428, 11'sd-558, 11'sd689}, {13'sd2320, 12'sd-1884, 13'sd-2753}, {10'sd-373, 13'sd-2331, 12'sd1249}},
{{12'sd-1222, 12'sd-1478, 10'sd329}, {12'sd-1447, 12'sd1538, 12'sd-1488}, {13'sd-2370, 13'sd2362, 12'sd1476}}},
{
{{12'sd1985, 12'sd-1532, 12'sd-1653}, {7'sd55, 12'sd-2003, 11'sd958}, {11'sd836, 12'sd-1803, 12'sd-1768}},
{{12'sd-1771, 12'sd1706, 12'sd-1639}, {12'sd-1988, 10'sd261, 12'sd-1343}, {12'sd-2047, 10'sd-452, 13'sd-2321}},
{{8'sd-114, 12'sd-2020, 10'sd261}, {13'sd-2631, 7'sd52, 12'sd1668}, {11'sd-549, 11'sd929, 13'sd2394}},
{{13'sd3223, 6'sd-16, 11'sd912}, {12'sd1497, 13'sd2539, 12'sd-1643}, {13'sd-3470, 7'sd-57, 13'sd-3504}},
{{12'sd-1513, 11'sd896, 11'sd-981}, {11'sd-531, 13'sd-2307, 9'sd235}, {11'sd-1023, 11'sd874, 12'sd1590}},
{{11'sd991, 9'sd199, 13'sd2435}, {13'sd2550, 11'sd725, 12'sd1715}, {12'sd1999, 11'sd-778, 12'sd1041}},
{{12'sd1632, 13'sd-2366, 10'sd326}, {12'sd1797, 12'sd-1378, 12'sd1506}, {12'sd-1382, 13'sd-3247, 11'sd-769}},
{{13'sd2100, 12'sd-1586, 12'sd1821}, {13'sd2466, 12'sd1062, 10'sd431}, {12'sd1056, 10'sd-293, 12'sd1254}},
{{13'sd-2177, 13'sd-2328, 13'sd-2444}, {12'sd1329, 12'sd1412, 12'sd1328}, {12'sd-1688, 11'sd-783, 13'sd-2763}},
{{11'sd-969, 12'sd1300, 13'sd-2325}, {13'sd-2459, 10'sd422, 13'sd2521}, {11'sd816, 12'sd1228, 12'sd1559}},
{{13'sd2391, 12'sd1759, 11'sd630}, {11'sd821, 9'sd161, 9'sd224}, {13'sd-2167, 13'sd-2497, 9'sd-208}},
{{11'sd-668, 9'sd-162, 12'sd1063}, {11'sd-1012, 11'sd-666, 12'sd1779}, {12'sd-1806, 9'sd170, 10'sd-347}},
{{7'sd43, 9'sd176, 12'sd1581}, {13'sd2363, 13'sd2832, 12'sd1983}, {6'sd26, 13'sd-3400, 11'sd-578}},
{{13'sd-2172, 12'sd-1988, 11'sd946}, {12'sd-1948, 12'sd-1897, 13'sd2563}, {13'sd-2684, 12'sd1250, 13'sd-2492}},
{{12'sd1707, 8'sd117, 11'sd-539}, {10'sd-336, 10'sd303, 12'sd1559}, {13'sd2604, 11'sd-692, 12'sd-2042}},
{{10'sd399, 12'sd1943, 11'sd-910}, {12'sd-1359, 12'sd-1484, 11'sd933}, {12'sd-1490, 12'sd1216, 13'sd2122}},
{{6'sd23, 9'sd253, 12'sd1227}, {11'sd926, 10'sd286, 11'sd869}, {12'sd-1916, 13'sd-2496, 12'sd-1163}},
{{13'sd-2740, 13'sd2722, 10'sd479}, {12'sd-1141, 10'sd328, 11'sd963}, {12'sd1030, 10'sd-333, 11'sd754}},
{{12'sd1857, 9'sd-175, 9'sd144}, {11'sd-544, 13'sd-2274, 12'sd-1726}, {13'sd-2148, 11'sd714, 12'sd-1275}},
{{13'sd2654, 12'sd-1568, 12'sd1680}, {12'sd-1978, 5'sd10, 11'sd-723}, {10'sd397, 13'sd2611, 8'sd-85}},
{{13'sd-2958, 11'sd-692, 10'sd-328}, {13'sd3437, 12'sd1877, 12'sd-1058}, {13'sd-2077, 12'sd-1236, 13'sd-2869}},
{{12'sd-1636, 12'sd2036, 10'sd-444}, {12'sd1512, 12'sd1916, 10'sd-287}, {11'sd-825, 10'sd-448, 12'sd-1228}},
{{13'sd-2218, 13'sd-2095, 12'sd-1877}, {12'sd1868, 11'sd964, 12'sd-1074}, {12'sd-1996, 12'sd-1845, 13'sd-2588}},
{{11'sd-658, 12'sd-2029, 11'sd514}, {11'sd707, 12'sd1650, 12'sd1125}, {13'sd-2200, 11'sd595, 12'sd1339}},
{{13'sd2587, 11'sd-862, 13'sd2086}, {9'sd180, 11'sd-728, 12'sd-1202}, {12'sd-1102, 12'sd1478, 13'sd-2373}},
{{10'sd-375, 11'sd1021, 12'sd1430}, {12'sd1657, 13'sd2620, 13'sd2482}, {12'sd-1213, 13'sd2662, 12'sd1923}},
{{12'sd1987, 12'sd-1460, 12'sd1688}, {13'sd-2630, 6'sd-20, 12'sd2012}, {8'sd-70, 13'sd2460, 13'sd-2119}},
{{11'sd815, 12'sd1031, 9'sd128}, {12'sd1679, 12'sd-2034, 12'sd2002}, {11'sd555, 10'sd304, 12'sd1727}},
{{13'sd2421, 11'sd-707, 12'sd-1835}, {10'sd372, 13'sd-2460, 11'sd-820}, {10'sd433, 13'sd-2415, 13'sd-2613}},
{{11'sd-870, 10'sd453, 13'sd2475}, {11'sd584, 13'sd2096, 12'sd1710}, {12'sd-1988, 11'sd-642, 9'sd161}},
{{12'sd1115, 12'sd-1447, 12'sd1704}, {11'sd522, 13'sd2712, 13'sd2261}, {10'sd-423, 12'sd-1207, 8'sd108}},
{{11'sd-889, 13'sd-2146, 11'sd738}, {12'sd-1655, 13'sd-2499, 10'sd349}, {12'sd1425, 13'sd-2074, 12'sd-1515}},
{{12'sd1190, 13'sd2068, 13'sd2373}, {13'sd-2098, 12'sd1871, 12'sd1145}, {9'sd-210, 13'sd2675, 12'sd1732}},
{{13'sd2725, 13'sd2415, 13'sd2345}, {12'sd-1086, 10'sd-350, 12'sd1167}, {6'sd-26, 10'sd267, 12'sd1468}},
{{13'sd-2619, 12'sd-1738, 10'sd-305}, {11'sd949, 10'sd349, 12'sd1306}, {12'sd-1903, 11'sd-1009, 12'sd1837}},
{{10'sd482, 13'sd2228, 13'sd-2253}, {13'sd2524, 12'sd1348, 12'sd1616}, {12'sd1125, 12'sd-1417, 13'sd-2410}},
{{11'sd570, 12'sd-1544, 13'sd2837}, {12'sd2044, 13'sd2480, 12'sd1660}, {13'sd-2624, 13'sd-2485, 13'sd2141}},
{{11'sd-825, 12'sd1389, 10'sd-281}, {11'sd-945, 13'sd2058, 12'sd-1312}, {11'sd832, 13'sd-2659, 12'sd-2005}},
{{13'sd-2076, 11'sd-687, 13'sd-2149}, {11'sd766, 9'sd-133, 10'sd-330}, {6'sd27, 11'sd852, 11'sd-1022}},
{{12'sd1719, 13'sd-2152, 12'sd1417}, {12'sd-1991, 12'sd1722, 12'sd1100}, {12'sd-1808, 12'sd-1974, 11'sd-1016}},
{{13'sd-3845, 9'sd-245, 10'sd508}, {13'sd-3300, 13'sd-2413, 11'sd550}, {13'sd-2702, 11'sd706, 11'sd-916}},
{{12'sd1112, 12'sd-2006, 11'sd950}, {13'sd-2554, 12'sd1769, 12'sd1525}, {12'sd1575, 13'sd2244, 12'sd-1166}},
{{11'sd631, 12'sd1549, 13'sd2172}, {12'sd-1031, 13'sd-2403, 12'sd-1345}, {12'sd1337, 12'sd1123, 12'sd-1673}},
{{11'sd552, 11'sd982, 13'sd2148}, {10'sd-469, 6'sd24, 11'sd904}, {13'sd2642, 11'sd844, 8'sd75}},
{{11'sd696, 9'sd-142, 12'sd-1751}, {8'sd-118, 12'sd-1723, 5'sd8}, {10'sd-312, 12'sd1363, 11'sd561}},
{{13'sd-2251, 13'sd2876, 11'sd552}, {12'sd1661, 12'sd-1737, 11'sd-525}, {12'sd-1191, 13'sd2383, 12'sd1664}},
{{11'sd-854, 10'sd-318, 10'sd-494}, {12'sd-1551, 12'sd-1334, 13'sd2340}, {11'sd-962, 13'sd2851, 11'sd983}},
{{13'sd-3081, 13'sd-2514, 13'sd-2417}, {11'sd-947, 12'sd1242, 11'sd-971}, {9'sd177, 13'sd-3776, 11'sd902}},
{{13'sd2173, 12'sd1957, 12'sd-1940}, {12'sd-1253, 12'sd1626, 12'sd1079}, {11'sd-625, 7'sd-47, 13'sd-3083}},
{{13'sd3562, 12'sd1090, 13'sd2726}, {10'sd488, 12'sd1719, 12'sd1218}, {14'sd4313, 12'sd1848, 10'sd501}},
{{10'sd-324, 12'sd1232, 12'sd1860}, {11'sd-701, 13'sd-2287, 11'sd-634}, {9'sd180, 11'sd999, 11'sd928}},
{{13'sd2562, 13'sd-2749, 12'sd1537}, {9'sd220, 11'sd-783, 13'sd2176}, {12'sd-1434, 12'sd1183, 11'sd876}},
{{9'sd-143, 12'sd1988, 12'sd1330}, {13'sd2294, 11'sd953, 10'sd351}, {12'sd-1179, 13'sd-2191, 9'sd-200}},
{{13'sd2640, 13'sd2739, 12'sd1472}, {13'sd2670, 12'sd-1451, 9'sd195}, {13'sd2786, 12'sd1420, 12'sd1055}},
{{13'sd-3716, 13'sd-3498, 13'sd-2759}, {12'sd-1710, 13'sd2825, 9'sd137}, {13'sd-2138, 12'sd-1803, 12'sd1045}},
{{7'sd-39, 12'sd1326, 9'sd-180}, {11'sd776, 11'sd544, 12'sd1650}, {12'sd1354, 11'sd-577, 12'sd1492}},
{{13'sd2636, 12'sd-1642, 11'sd-827}, {10'sd-291, 12'sd-1574, 7'sd38}, {13'sd-2722, 12'sd1985, 12'sd-1376}},
{{11'sd610, 11'sd784, 13'sd-2399}, {13'sd2538, 12'sd-1049, 10'sd488}, {13'sd2799, 12'sd-1798, 12'sd-1185}},
{{12'sd1471, 13'sd2752, 12'sd-2013}, {11'sd794, 11'sd673, 12'sd-1263}, {11'sd-756, 12'sd-1117, 13'sd2329}},
{{12'sd-1211, 12'sd-1096, 11'sd937}, {11'sd512, 10'sd292, 11'sd-941}, {10'sd-428, 11'sd985, 12'sd-1385}},
{{12'sd1162, 11'sd685, 12'sd1197}, {11'sd986, 12'sd-1130, 11'sd1010}, {13'sd2765, 12'sd1194, 11'sd-932}},
{{13'sd2154, 13'sd3003, 13'sd2129}, {12'sd-2019, 12'sd1256, 10'sd-438}, {13'sd-2179, 11'sd646, 12'sd-1040}},
{{12'sd1820, 13'sd2718, 12'sd-1384}, {11'sd727, 12'sd-1770, 13'sd2448}, {12'sd1727, 10'sd-441, 12'sd1055}},
{{11'sd513, 12'sd-1318, 12'sd-1917}, {13'sd-2399, 12'sd-1095, 12'sd1485}, {12'sd-1930, 12'sd1565, 13'sd2740}}},
{
{{11'sd-733, 12'sd1471, 12'sd-1032}, {13'sd2450, 10'sd-409, 12'sd1574}, {11'sd-868, 12'sd1993, 12'sd1258}},
{{12'sd-1692, 9'sd-180, 11'sd886}, {12'sd1637, 12'sd-2014, 11'sd-532}, {12'sd-1831, 10'sd371, 8'sd90}},
{{13'sd-2275, 12'sd1877, 8'sd-117}, {12'sd1598, 9'sd250, 13'sd-2159}, {12'sd-1069, 13'sd-2225, 12'sd-1454}},
{{13'sd-2317, 11'sd543, 13'sd2229}, {12'sd1911, 12'sd-1048, 12'sd1165}, {9'sd141, 11'sd802, 11'sd651}},
{{9'sd134, 12'sd-1709, 13'sd2542}, {11'sd716, 12'sd1815, 13'sd-2650}, {12'sd-1561, 9'sd210, 12'sd-1881}},
{{13'sd2108, 13'sd2176, 12'sd1508}, {11'sd-643, 13'sd2639, 12'sd1058}, {10'sd-318, 11'sd-749, 13'sd2425}},
{{12'sd-1925, 12'sd1172, 12'sd-1711}, {12'sd1528, 12'sd-1478, 12'sd-1748}, {12'sd-1161, 12'sd1308, 13'sd3069}},
{{12'sd-1068, 11'sd687, 13'sd-3289}, {12'sd1088, 11'sd-914, 13'sd-2480}, {12'sd-1998, 12'sd-1261, 10'sd-345}},
{{11'sd-595, 13'sd3100, 13'sd2687}, {11'sd-887, 13'sd2890, 11'sd-552}, {12'sd-1164, 13'sd-2402, 13'sd-2749}},
{{13'sd2421, 11'sd738, 12'sd1697}, {10'sd-286, 13'sd2606, 9'sd-148}, {13'sd2356, 12'sd-1400, 9'sd-211}},
{{12'sd1326, 13'sd-2741, 13'sd-2765}, {12'sd1691, 13'sd-2955, 11'sd-904}, {9'sd-135, 12'sd1811, 12'sd-1599}},
{{13'sd-3164, 12'sd-1759, 13'sd-2617}, {12'sd1801, 11'sd-971, 12'sd1654}, {13'sd-2545, 13'sd-2098, 11'sd616}},
{{10'sd277, 11'sd-773, 13'sd-2205}, {12'sd-1433, 11'sd739, 13'sd2072}, {13'sd3647, 13'sd2863, 9'sd170}},
{{13'sd-2926, 12'sd-1520, 11'sd969}, {13'sd2432, 12'sd-1663, 11'sd839}, {12'sd-1650, 13'sd2611, 12'sd-1521}},
{{12'sd-1774, 7'sd61, 12'sd-1642}, {11'sd-963, 11'sd-657, 12'sd-1977}, {13'sd-2809, 9'sd-236, 7'sd35}},
{{12'sd1493, 12'sd-2012, 12'sd1965}, {11'sd787, 10'sd-271, 11'sd555}, {11'sd-562, 13'sd2270, 12'sd1069}},
{{12'sd1917, 13'sd2852, 11'sd641}, {11'sd-636, 13'sd2811, 13'sd2207}, {13'sd2235, 11'sd-816, 11'sd795}},
{{12'sd1905, 11'sd-701, 11'sd-666}, {12'sd1976, 13'sd-2522, 9'sd-146}, {13'sd2853, 11'sd-542, 11'sd-914}},
{{13'sd-2615, 11'sd-670, 8'sd72}, {11'sd754, 11'sd766, 12'sd1822}, {11'sd528, 13'sd-2187, 12'sd-1969}},
{{11'sd843, 12'sd1186, 13'sd-2519}, {11'sd-541, 12'sd-1510, 9'sd-174}, {12'sd-1196, 13'sd-2145, 13'sd-2555}},
{{11'sd673, 11'sd850, 9'sd188}, {13'sd2899, 13'sd-2276, 13'sd2953}, {9'sd192, 11'sd-1014, 9'sd-172}},
{{10'sd333, 12'sd1075, 13'sd-2858}, {12'sd1502, 9'sd197, 12'sd2004}, {13'sd2311, 13'sd2240, 13'sd-2424}},
{{12'sd-1573, 9'sd-206, 10'sd-472}, {12'sd1658, 12'sd-1712, 11'sd-893}, {12'sd-1051, 10'sd285, 13'sd-2419}},
{{13'sd2172, 12'sd1547, 12'sd-1634}, {13'sd-2169, 12'sd-1767, 11'sd-685}, {10'sd440, 11'sd-656, 11'sd597}},
{{13'sd-2371, 11'sd579, 13'sd-2717}, {12'sd-1472, 13'sd-2145, 11'sd733}, {13'sd-2961, 13'sd-2894, 12'sd-1076}},
{{12'sd-1793, 11'sd908, 12'sd-1917}, {13'sd2214, 11'sd901, 11'sd703}, {12'sd1339, 12'sd1345, 13'sd-2096}},
{{13'sd3030, 12'sd1040, 12'sd1778}, {11'sd888, 9'sd217, 11'sd-672}, {13'sd2503, 12'sd-1767, 12'sd-1336}},
{{13'sd-2462, 9'sd239, 10'sd-397}, {12'sd-1514, 8'sd86, 12'sd-1938}, {9'sd233, 12'sd-1873, 11'sd819}},
{{12'sd-1097, 12'sd1469, 8'sd-121}, {12'sd-1388, 12'sd1929, 13'sd2839}, {12'sd1414, 11'sd606, 7'sd-48}},
{{13'sd2291, 9'sd191, 11'sd547}, {12'sd1668, 10'sd453, 13'sd-2760}, {13'sd-2825, 11'sd-985, 12'sd-1994}},
{{12'sd-1107, 13'sd-3054, 13'sd-2318}, {12'sd1118, 11'sd559, 13'sd-2363}, {13'sd2685, 12'sd1706, 12'sd-1318}},
{{10'sd-315, 9'sd200, 11'sd851}, {13'sd2784, 12'sd1826, 13'sd2361}, {12'sd-1852, 12'sd1198, 12'sd-1064}},
{{13'sd-3320, 13'sd-2928, 12'sd2027}, {12'sd-1718, 9'sd182, 12'sd-1257}, {13'sd2683, 11'sd-605, 12'sd1963}},
{{12'sd-1507, 12'sd-1467, 9'sd-242}, {12'sd-1693, 13'sd-2898, 11'sd774}, {12'sd-1053, 11'sd-627, 12'sd-1844}},
{{11'sd-944, 13'sd2116, 11'sd801}, {12'sd-1310, 12'sd1957, 12'sd1256}, {13'sd2146, 11'sd1003, 9'sd-158}},
{{13'sd-2575, 12'sd-2017, 12'sd1462}, {12'sd-1242, 5'sd-8, 12'sd-1769}, {13'sd2192, 11'sd-748, 10'sd-267}},
{{13'sd2532, 13'sd2244, 12'sd-1214}, {11'sd-1012, 13'sd-2203, 12'sd1945}, {12'sd1807, 13'sd3021, 10'sd-399}},
{{9'sd-234, 8'sd127, 9'sd176}, {9'sd-249, 12'sd-1746, 13'sd-2397}, {10'sd342, 12'sd1691, 12'sd1600}},
{{13'sd3015, 12'sd1352, 13'sd2933}, {13'sd-2408, 13'sd-2265, 11'sd-641}, {10'sd-331, 12'sd-1972, 13'sd2379}},
{{12'sd-1141, 10'sd501, 12'sd-2025}, {11'sd-550, 12'sd1824, 10'sd-446}, {12'sd1450, 12'sd1359, 12'sd-1519}},
{{13'sd-2370, 12'sd-1787, 13'sd-2453}, {12'sd1566, 12'sd1707, 12'sd1867}, {13'sd2604, 12'sd-1316, 12'sd-1076}},
{{12'sd-1164, 10'sd457, 12'sd-1507}, {11'sd-811, 11'sd-928, 12'sd2035}, {11'sd875, 12'sd1191, 13'sd3231}},
{{12'sd-1035, 13'sd-2391, 11'sd-783}, {11'sd891, 12'sd1833, 13'sd3015}, {11'sd-962, 11'sd738, 13'sd2216}},
{{11'sd-642, 7'sd55, 10'sd-299}, {12'sd-1479, 11'sd772, 11'sd-1018}, {13'sd2387, 13'sd-2540, 11'sd-819}},
{{12'sd1998, 12'sd1592, 12'sd1596}, {12'sd-1323, 13'sd2917, 9'sd-150}, {13'sd2244, 11'sd785, 11'sd-869}},
{{13'sd-2361, 13'sd2285, 12'sd-1159}, {10'sd274, 12'sd2027, 12'sd1793}, {13'sd-2509, 10'sd390, 11'sd-833}},
{{12'sd1292, 11'sd-845, 11'sd-904}, {12'sd1336, 12'sd-1591, 10'sd-313}, {13'sd2135, 10'sd336, 13'sd-2334}},
{{12'sd-1325, 13'sd2295, 10'sd288}, {13'sd-2197, 10'sd-432, 11'sd-550}, {13'sd2224, 13'sd2759, 13'sd3277}},
{{13'sd3022, 9'sd-169, 10'sd-389}, {12'sd1671, 13'sd-2559, 12'sd-1358}, {12'sd-1271, 13'sd-2316, 12'sd-1758}},
{{8'sd106, 13'sd2972, 7'sd-46}, {13'sd-2356, 13'sd-3044, 10'sd-455}, {13'sd-2298, 13'sd-2955, 12'sd1134}},
{{12'sd-1421, 12'sd-1285, 12'sd-1367}, {13'sd-3517, 10'sd-317, 11'sd630}, {13'sd-2486, 11'sd-968, 11'sd742}},
{{12'sd-1248, 13'sd2520, 12'sd-1823}, {12'sd-1952, 10'sd487, 11'sd584}, {10'sd403, 12'sd-1037, 9'sd-204}},
{{11'sd666, 8'sd-108, 6'sd-29}, {12'sd1582, 13'sd2486, 13'sd2177}, {12'sd1409, 11'sd-772, 12'sd1217}},
{{8'sd112, 10'sd-372, 6'sd29}, {12'sd-1105, 12'sd-1554, 10'sd494}, {12'sd-1690, 12'sd1536, 13'sd2468}},
{{12'sd1691, 12'sd1111, 13'sd2119}, {12'sd-1113, 12'sd1252, 12'sd-1692}, {13'sd2220, 12'sd1248, 12'sd1538}},
{{12'sd-1717, 13'sd-2399, 12'sd1682}, {12'sd-1450, 13'sd-2091, 13'sd-2481}, {12'sd1588, 10'sd-347, 13'sd2676}},
{{13'sd-2848, 13'sd2318, 12'sd-1897}, {12'sd-1233, 13'sd2463, 12'sd1515}, {11'sd766, 9'sd247, 9'sd-241}},
{{11'sd548, 13'sd2476, 13'sd-2666}, {7'sd48, 11'sd-614, 9'sd229}, {11'sd708, 13'sd2099, 13'sd-2243}},
{{12'sd-1797, 11'sd-711, 10'sd326}, {13'sd2484, 8'sd-103, 12'sd1149}, {9'sd-253, 13'sd3013, 11'sd-854}},
{{12'sd-1529, 12'sd1365, 12'sd1077}, {12'sd-1664, 11'sd680, 12'sd-1697}, {12'sd-1215, 7'sd-52, 5'sd-11}},
{{12'sd1050, 12'sd-1041, 13'sd2423}, {13'sd2377, 13'sd2312, 8'sd-81}, {12'sd-1909, 13'sd-2352, 12'sd-1754}},
{{13'sd-2203, 13'sd-2357, 12'sd1236}, {13'sd-2389, 7'sd55, 13'sd-2597}, {12'sd-1055, 9'sd-221, 12'sd-1338}},
{{8'sd92, 13'sd-2898, 11'sd673}, {13'sd2226, 12'sd1735, 12'sd2012}, {12'sd1603, 11'sd686, 12'sd-1922}},
{{13'sd-2208, 12'sd1401, 9'sd-178}, {11'sd-1001, 10'sd-449, 12'sd1528}, {10'sd435, 11'sd-632, 12'sd-1614}}},
{
{{13'sd2281, 10'sd415, 11'sd-581}, {13'sd-2939, 12'sd1832, 12'sd-1083}, {7'sd41, 9'sd-215, 12'sd-1447}},
{{12'sd-1662, 13'sd2194, 12'sd1089}, {11'sd655, 11'sd-566, 13'sd-2875}, {12'sd1169, 8'sd72, 11'sd847}},
{{13'sd3157, 13'sd3204, 12'sd1975}, {13'sd2606, 13'sd2333, 9'sd-248}, {13'sd-2550, 13'sd2187, 12'sd-1192}},
{{11'sd-926, 12'sd-1422, 12'sd-1685}, {10'sd356, 12'sd1913, 9'sd-145}, {12'sd1434, 12'sd1969, 13'sd-3265}},
{{13'sd2607, 12'sd1741, 12'sd-1459}, {9'sd-138, 12'sd2014, 13'sd2617}, {13'sd2078, 7'sd-48, 13'sd-2398}},
{{10'sd296, 12'sd1232, 11'sd807}, {12'sd1312, 12'sd1387, 13'sd2281}, {11'sd-843, 11'sd575, 12'sd-1769}},
{{11'sd652, 9'sd176, 12'sd-1821}, {12'sd-1197, 12'sd-1907, 11'sd-684}, {13'sd3459, 12'sd-1165, 13'sd2076}},
{{12'sd1473, 11'sd713, 11'sd-680}, {11'sd862, 12'sd1214, 11'sd-632}, {12'sd-1429, 12'sd-1406, 11'sd-525}},
{{12'sd-1486, 12'sd1037, 13'sd2598}, {11'sd-594, 10'sd402, 12'sd-1726}, {10'sd-317, 13'sd-2453, 9'sd134}},
{{12'sd1179, 12'sd-1096, 12'sd1929}, {12'sd1633, 12'sd-1403, 13'sd2408}, {10'sd342, 11'sd-560, 12'sd-1184}},
{{13'sd-2640, 13'sd2079, 12'sd-1319}, {11'sd-926, 11'sd807, 9'sd-142}, {13'sd-2463, 12'sd1185, 11'sd517}},
{{11'sd-574, 11'sd-517, 10'sd-368}, {11'sd-556, 11'sd-976, 11'sd775}, {13'sd2233, 12'sd-1491, 11'sd673}},
{{13'sd-3135, 12'sd-1404, 12'sd1574}, {13'sd-3213, 13'sd-2362, 11'sd-908}, {12'sd1447, 11'sd-653, 12'sd-1137}},
{{12'sd-1652, 12'sd1315, 13'sd-2214}, {11'sd-718, 11'sd-545, 8'sd104}, {12'sd-1649, 13'sd2553, 10'sd-396}},
{{11'sd-952, 12'sd1675, 12'sd-1274}, {12'sd-1327, 10'sd-495, 10'sd366}, {13'sd-2809, 11'sd713, 12'sd1657}},
{{7'sd-61, 13'sd-2457, 11'sd726}, {12'sd1797, 11'sd690, 13'sd2645}, {13'sd-2323, 11'sd-585, 13'sd2150}},
{{10'sd-456, 13'sd2699, 13'sd2722}, {11'sd-700, 13'sd2148, 11'sd781}, {13'sd-2210, 13'sd2387, 12'sd1375}},
{{12'sd1899, 13'sd-3185, 11'sd843}, {12'sd-1127, 10'sd-480, 12'sd1964}, {9'sd-149, 11'sd977, 13'sd-2120}},
{{12'sd-1259, 8'sd-97, 11'sd-857}, {12'sd1716, 12'sd1815, 12'sd1918}, {13'sd2642, 11'sd-657, 12'sd1343}},
{{12'sd-1762, 12'sd-1308, 11'sd-702}, {12'sd-1900, 12'sd1332, 12'sd-1129}, {12'sd-1440, 10'sd326, 12'sd-1257}},
{{13'sd2792, 10'sd-393, 13'sd-2862}, {12'sd1519, 6'sd-24, 12'sd-1155}, {9'sd211, 12'sd2009, 12'sd-1542}},
{{11'sd532, 12'sd-1797, 12'sd1942}, {10'sd-471, 12'sd1355, 12'sd-1755}, {11'sd-641, 13'sd2525, 11'sd705}},
{{9'sd140, 12'sd1774, 13'sd2220}, {9'sd-206, 11'sd-956, 12'sd1688}, {13'sd2052, 12'sd1183, 13'sd-2426}},
{{13'sd-2382, 13'sd2215, 13'sd-2775}, {10'sd-305, 11'sd-819, 13'sd-2444}, {12'sd1751, 12'sd-1563, 9'sd-213}},
{{13'sd2346, 12'sd-1285, 11'sd1014}, {12'sd-1748, 12'sd-1935, 13'sd2769}, {12'sd1454, 11'sd-981, 10'sd-342}},
{{12'sd1611, 10'sd294, 12'sd-1300}, {12'sd1202, 13'sd-2443, 11'sd-692}, {11'sd-605, 12'sd-1622, 12'sd-1623}},
{{13'sd2347, 10'sd-472, 13'sd-2410}, {13'sd-2133, 11'sd-866, 11'sd662}, {11'sd884, 10'sd-364, 13'sd-2670}},
{{12'sd-1463, 11'sd-785, 12'sd-1860}, {12'sd-1880, 13'sd2631, 11'sd-745}, {13'sd2569, 12'sd-1916, 12'sd-1889}},
{{12'sd1288, 13'sd-2125, 12'sd1116}, {7'sd-32, 10'sd369, 9'sd135}, {10'sd-338, 12'sd1980, 10'sd439}},
{{10'sd323, 11'sd-964, 13'sd2489}, {13'sd-2312, 8'sd123, 12'sd1123}, {12'sd-1082, 12'sd1155, 12'sd-1700}},
{{12'sd-2041, 8'sd-106, 13'sd-3904}, {11'sd-567, 12'sd1195, 12'sd1264}, {8'sd116, 13'sd3070, 10'sd415}},
{{12'sd-1336, 12'sd1479, 7'sd37}, {11'sd-522, 11'sd730, 12'sd-1916}, {11'sd-671, 12'sd1280, 11'sd889}},
{{12'sd-1580, 10'sd-480, 10'sd496}, {12'sd-1887, 12'sd-1608, 12'sd1145}, {10'sd459, 11'sd1015, 12'sd-1138}},
{{13'sd2348, 13'sd2520, 12'sd-1671}, {11'sd518, 9'sd-134, 13'sd-2405}, {9'sd-253, 10'sd-510, 12'sd1462}},
{{11'sd965, 13'sd2460, 12'sd1075}, {12'sd1284, 12'sd-1750, 12'sd1041}, {12'sd1635, 12'sd1624, 13'sd2817}},
{{13'sd-2871, 11'sd891, 13'sd-2058}, {12'sd-1133, 12'sd1489, 12'sd1325}, {10'sd376, 7'sd33, 13'sd-2361}},
{{10'sd404, 12'sd-1169, 12'sd1794}, {10'sd351, 11'sd-667, 13'sd-2391}, {12'sd1356, 12'sd-1831, 11'sd959}},
{{12'sd1065, 12'sd1513, 11'sd-884}, {12'sd1764, 11'sd930, 12'sd-1154}, {13'sd2581, 11'sd-678, 12'sd-1740}},
{{10'sd-366, 12'sd-1250, 12'sd1643}, {13'sd-2858, 11'sd1019, 11'sd-907}, {13'sd-2292, 13'sd-2351, 12'sd-1275}},
{{13'sd-2325, 8'sd-68, 12'sd1808}, {12'sd1928, 12'sd-1741, 12'sd-1130}, {13'sd-3030, 13'sd-3416, 13'sd-3078}},
{{7'sd-38, 12'sd1847, 11'sd594}, {9'sd-147, 9'sd-146, 13'sd-2532}, {11'sd-661, 12'sd-1119, 12'sd1921}},
{{13'sd3028, 8'sd-68, 13'sd2399}, {13'sd-3496, 12'sd-1255, 12'sd1877}, {9'sd216, 13'sd2403, 12'sd1063}},
{{12'sd-1070, 13'sd-2423, 11'sd519}, {10'sd439, 13'sd-2997, 12'sd-1441}, {12'sd1948, 11'sd881, 12'sd1678}},
{{12'sd1615, 13'sd-2194, 13'sd-2228}, {12'sd1148, 7'sd45, 11'sd-537}, {12'sd-1576, 11'sd-1002, 12'sd-1420}},
{{11'sd725, 10'sd-379, 13'sd2823}, {12'sd-1899, 12'sd1465, 12'sd1348}, {7'sd-37, 13'sd2131, 12'sd-1852}},
{{8'sd-108, 13'sd-2135, 13'sd-2382}, {13'sd2497, 11'sd950, 11'sd631}, {11'sd-903, 9'sd145, 12'sd2032}},
{{12'sd-1513, 11'sd666, 13'sd2244}, {13'sd-2694, 13'sd-2480, 10'sd458}, {9'sd194, 10'sd-330, 11'sd-801}},
{{13'sd2872, 6'sd30, 10'sd321}, {12'sd-1100, 13'sd-2529, 12'sd-1062}, {10'sd-326, 8'sd68, 9'sd-242}},
{{11'sd-571, 12'sd-1640, 13'sd-2067}, {13'sd2845, 13'sd3084, 12'sd1618}, {11'sd-825, 11'sd-965, 12'sd-2011}},
{{11'sd569, 11'sd-588, 11'sd1011}, {13'sd3075, 13'sd2574, 13'sd2153}, {13'sd3208, 12'sd-1608, 12'sd-1685}},
{{9'sd206, 13'sd2301, 12'sd2010}, {13'sd-2332, 11'sd-701, 11'sd-731}, {13'sd-3016, 12'sd1700, 9'sd167}},
{{11'sd-991, 12'sd-1889, 10'sd453}, {12'sd1095, 12'sd1992, 13'sd-2795}, {12'sd-1204, 10'sd-379, 13'sd2314}},
{{5'sd-15, 13'sd-2246, 12'sd1290}, {10'sd-456, 7'sd48, 12'sd-1489}, {13'sd2142, 13'sd2474, 13'sd-2742}},
{{13'sd2324, 12'sd-1959, 12'sd1075}, {12'sd-1440, 9'sd187, 6'sd-30}, {13'sd-2407, 13'sd-2568, 11'sd549}},
{{11'sd-708, 13'sd2061, 11'sd-799}, {12'sd-1698, 13'sd-2846, 12'sd-1441}, {13'sd-3071, 12'sd1746, 13'sd3427}},
{{13'sd2726, 11'sd1008, 10'sd-265}, {13'sd-2290, 12'sd-1674, 12'sd1452}, {12'sd1573, 13'sd-2127, 13'sd2527}},
{{13'sd-2313, 13'sd-2086, 10'sd449}, {12'sd-1310, 13'sd-2596, 12'sd-1516}, {13'sd-2423, 11'sd800, 13'sd-2246}},
{{11'sd-602, 10'sd-448, 11'sd727}, {12'sd1611, 11'sd-525, 12'sd-1702}, {8'sd-95, 12'sd1530, 11'sd-645}},
{{11'sd823, 10'sd-488, 12'sd1087}, {10'sd460, 13'sd-3234, 12'sd-1284}, {12'sd1131, 13'sd2607, 11'sd-970}},
{{13'sd-2620, 12'sd-1534, 13'sd2091}, {10'sd489, 12'sd1035, 12'sd2000}, {10'sd-378, 10'sd-417, 10'sd372}},
{{12'sd1093, 13'sd2502, 9'sd242}, {11'sd908, 13'sd2710, 11'sd-973}, {11'sd-597, 9'sd214, 11'sd681}},
{{10'sd-500, 12'sd1609, 7'sd-42}, {11'sd599, 12'sd-1455, 13'sd-3238}, {12'sd-1133, 12'sd-1327, 10'sd476}},
{{11'sd-667, 12'sd1632, 9'sd253}, {13'sd-2254, 12'sd1169, 10'sd382}, {10'sd393, 13'sd-2149, 12'sd1603}},
{{10'sd386, 13'sd2287, 11'sd-813}, {12'sd1914, 13'sd2820, 12'sd-1067}, {11'sd738, 13'sd2251, 11'sd-982}}},
{
{{13'sd2487, 13'sd2417, 10'sd-353}, {11'sd626, 11'sd686, 13'sd2452}, {12'sd1678, 12'sd1221, 7'sd-50}},
{{11'sd-855, 10'sd-438, 8'sd77}, {9'sd-181, 11'sd-724, 13'sd2271}, {12'sd-1478, 13'sd2198, 11'sd-578}},
{{12'sd1607, 12'sd1259, 13'sd2754}, {12'sd1389, 13'sd-2271, 13'sd-2463}, {13'sd-2162, 12'sd-1579, 13'sd2067}},
{{12'sd-2004, 13'sd-2896, 11'sd839}, {8'sd115, 9'sd-243, 10'sd332}, {13'sd-2148, 11'sd-777, 13'sd-2680}},
{{12'sd1834, 13'sd2973, 12'sd-1173}, {13'sd2165, 13'sd-2129, 9'sd-194}, {11'sd-1022, 13'sd2852, 13'sd2490}},
{{11'sd557, 11'sd690, 12'sd-1127}, {11'sd-637, 13'sd2178, 11'sd647}, {9'sd-185, 9'sd-183, 13'sd2424}},
{{12'sd-1553, 12'sd1331, 13'sd-2744}, {12'sd1956, 11'sd-885, 12'sd1314}, {13'sd2121, 9'sd-241, 12'sd-1189}},
{{12'sd-1321, 13'sd2068, 12'sd1721}, {12'sd1783, 10'sd405, 12'sd1973}, {11'sd634, 12'sd1489, 11'sd-524}},
{{10'sd494, 12'sd-1282, 13'sd-2665}, {12'sd1143, 13'sd-3103, 12'sd1629}, {12'sd1136, 10'sd-407, 12'sd-1331}},
{{11'sd671, 11'sd799, 12'sd1939}, {11'sd1003, 6'sd-27, 12'sd1570}, {12'sd1709, 11'sd-695, 13'sd-2322}},
{{11'sd929, 13'sd-3283, 10'sd504}, {13'sd-3116, 13'sd-2499, 13'sd-2849}, {10'sd413, 12'sd-1414, 12'sd1224}},
{{11'sd989, 13'sd2189, 12'sd-1062}, {11'sd-845, 13'sd-2143, 13'sd2155}, {12'sd-1528, 12'sd-1108, 11'sd-981}},
{{13'sd-2531, 11'sd-722, 13'sd-3230}, {12'sd-1834, 12'sd-1212, 11'sd-898}, {13'sd2054, 10'sd307, 12'sd-1354}},
{{10'sd310, 13'sd2416, 13'sd2324}, {12'sd-1939, 11'sd631, 11'sd-834}, {11'sd-639, 12'sd-1710, 12'sd1468}},
{{6'sd-17, 12'sd1168, 8'sd-114}, {12'sd-1846, 13'sd2233, 11'sd-807}, {11'sd583, 13'sd-2228, 10'sd437}},
{{11'sd622, 13'sd2237, 12'sd-1145}, {11'sd739, 12'sd1336, 11'sd-654}, {12'sd-1245, 11'sd-752, 11'sd-975}},
{{12'sd1331, 12'sd1725, 13'sd2147}, {9'sd-166, 12'sd1437, 13'sd2328}, {11'sd-681, 13'sd-2130, 11'sd740}},
{{13'sd2998, 10'sd318, 11'sd-843}, {13'sd2366, 10'sd399, 12'sd-1890}, {11'sd660, 12'sd1610, 12'sd1484}},
{{12'sd1516, 12'sd-1644, 13'sd2456}, {13'sd2460, 13'sd2480, 13'sd2466}, {6'sd28, 10'sd281, 12'sd-1166}},
{{10'sd-479, 13'sd-2799, 12'sd1202}, {13'sd-2693, 11'sd939, 11'sd529}, {12'sd-1405, 11'sd908, 12'sd1357}},
{{12'sd-1677, 12'sd1236, 10'sd455}, {13'sd-2229, 12'sd1474, 10'sd396}, {11'sd951, 12'sd-1518, 13'sd2516}},
{{12'sd-1693, 13'sd-3541, 13'sd-2628}, {12'sd-1367, 13'sd-3089, 8'sd-94}, {13'sd-2757, 13'sd-2763, 13'sd-2874}},
{{12'sd1111, 11'sd974, 12'sd2020}, {12'sd1141, 11'sd-568, 7'sd52}, {13'sd-2515, 12'sd1297, 7'sd61}},
{{12'sd-1159, 12'sd1611, 13'sd2303}, {12'sd1122, 10'sd313, 12'sd-2034}, {12'sd1135, 12'sd-1466, 12'sd-1156}},
{{11'sd-980, 12'sd1092, 11'sd-843}, {12'sd-1032, 12'sd-1091, 12'sd1544}, {13'sd-2997, 12'sd1829, 11'sd-873}},
{{9'sd-201, 12'sd-1924, 12'sd1927}, {12'sd1156, 12'sd1159, 11'sd-645}, {13'sd-2438, 12'sd-1794, 12'sd-1156}},
{{9'sd-135, 13'sd2380, 11'sd-704}, {11'sd-717, 11'sd964, 12'sd-1218}, {9'sd193, 13'sd2979, 10'sd-488}},
{{13'sd-2784, 10'sd-511, 13'sd-2363}, {12'sd-1196, 11'sd-981, 12'sd-1072}, {10'sd349, 11'sd996, 12'sd1688}},
{{12'sd-1128, 12'sd1730, 12'sd1953}, {10'sd-375, 10'sd420, 13'sd-2279}, {12'sd-2042, 12'sd-1687, 11'sd890}},
{{12'sd-1820, 12'sd1835, 12'sd1906}, {13'sd-2086, 12'sd1075, 13'sd2458}, {13'sd-2541, 10'sd-448, 10'sd-390}},
{{13'sd2125, 13'sd2625, 12'sd1976}, {13'sd2905, 11'sd-915, 12'sd-1876}, {13'sd2082, 13'sd3720, 11'sd-771}},
{{10'sd316, 13'sd2465, 13'sd-2069}, {11'sd-913, 6'sd30, 13'sd2853}, {13'sd-2256, 11'sd-772, 12'sd-1563}},
{{12'sd-1390, 12'sd-1288, 12'sd1244}, {12'sd-1788, 12'sd1248, 11'sd-779}, {11'sd-907, 12'sd-2034, 9'sd170}},
{{12'sd-1329, 12'sd-1686, 13'sd-2276}, {9'sd-237, 12'sd1776, 12'sd-1544}, {12'sd-1678, 12'sd1877, 10'sd432}},
{{11'sd-556, 12'sd1294, 12'sd-1528}, {12'sd-1859, 12'sd1721, 11'sd-837}, {12'sd1427, 13'sd2486, 12'sd-1537}},
{{12'sd-1519, 12'sd-1546, 11'sd-792}, {11'sd914, 11'sd866, 12'sd1208}, {12'sd-1297, 13'sd-2726, 10'sd470}},
{{12'sd-1655, 11'sd-868, 9'sd-145}, {12'sd-1639, 11'sd-780, 11'sd1007}, {12'sd-1922, 11'sd-741, 12'sd1297}},
{{12'sd-1101, 12'sd-2040, 12'sd1332}, {12'sd-1265, 13'sd2053, 13'sd2276}, {7'sd-43, 10'sd459, 10'sd468}},
{{10'sd475, 13'sd2158, 11'sd-721}, {10'sd452, 11'sd669, 13'sd2795}, {10'sd-371, 13'sd2880, 13'sd2469}},
{{10'sd388, 12'sd1300, 12'sd1407}, {11'sd-974, 11'sd-725, 8'sd73}, {9'sd195, 9'sd-222, 12'sd-1865}},
{{12'sd1403, 8'sd99, 13'sd-2789}, {13'sd2522, 9'sd245, 13'sd-2482}, {12'sd-1553, 13'sd2161, 12'sd1666}},
{{13'sd-2780, 13'sd2501, 12'sd1333}, {13'sd2104, 13'sd2473, 11'sd805}, {13'sd-3202, 13'sd2317, 12'sd1736}},
{{12'sd1705, 8'sd-80, 11'sd996}, {12'sd1176, 12'sd-1582, 13'sd2764}, {8'sd-126, 10'sd381, 12'sd1905}},
{{11'sd-586, 12'sd1699, 12'sd1220}, {12'sd1584, 12'sd1387, 11'sd-729}, {12'sd2038, 11'sd-1015, 12'sd-1412}},
{{12'sd-1543, 12'sd1663, 9'sd145}, {11'sd1007, 10'sd473, 12'sd1393}, {12'sd-1831, 11'sd-591, 13'sd2303}},
{{11'sd-744, 12'sd-1453, 13'sd-2975}, {13'sd-2711, 12'sd-2026, 13'sd-2263}, {12'sd1092, 10'sd292, 12'sd-1444}},
{{13'sd-2881, 9'sd184, 12'sd-1346}, {13'sd-3147, 13'sd-2105, 12'sd-1683}, {12'sd-1654, 12'sd-1805, 13'sd-2184}},
{{13'sd-2340, 13'sd2394, 13'sd2329}, {12'sd1443, 13'sd-2417, 6'sd-25}, {10'sd479, 11'sd-995, 13'sd-2553}},
{{13'sd2170, 8'sd-92, 11'sd-841}, {12'sd1298, 10'sd266, 13'sd-2262}, {11'sd-897, 11'sd710, 12'sd1397}},
{{12'sd-1114, 11'sd-805, 13'sd3197}, {11'sd-574, 11'sd-905, 12'sd-1589}, {12'sd1160, 12'sd1584, 13'sd-2361}},
{{12'sd-1859, 11'sd773, 11'sd-998}, {13'sd2608, 13'sd2512, 12'sd1969}, {11'sd-846, 12'sd1519, 13'sd3519}},
{{10'sd-299, 11'sd-839, 12'sd-1214}, {13'sd2589, 13'sd-2311, 12'sd1782}, {11'sd676, 12'sd-1192, 12'sd-1198}},
{{13'sd-2789, 12'sd-1414, 11'sd-606}, {12'sd-1304, 13'sd2428, 12'sd-1349}, {11'sd-915, 11'sd991, 10'sd-466}},
{{10'sd296, 9'sd141, 11'sd868}, {12'sd-1169, 9'sd189, 12'sd-1712}, {13'sd2773, 12'sd-1594, 10'sd269}},
{{13'sd-2725, 9'sd198, 10'sd482}, {11'sd645, 10'sd-437, 12'sd1733}, {11'sd980, 12'sd1074, 13'sd2314}},
{{11'sd-740, 7'sd-49, 12'sd-1129}, {6'sd-20, 13'sd-2924, 12'sd-1241}, {12'sd1079, 11'sd658, 12'sd-1187}},
{{12'sd1966, 13'sd-2213, 10'sd500}, {12'sd-1672, 12'sd1798, 12'sd-1234}, {12'sd-1150, 12'sd1951, 13'sd2496}},
{{13'sd2766, 13'sd-2338, 13'sd2071}, {12'sd-1580, 8'sd-125, 13'sd2233}, {13'sd2500, 13'sd-2737, 12'sd1669}},
{{13'sd-2540, 12'sd1253, 10'sd-382}, {8'sd-124, 10'sd-298, 13'sd2351}, {10'sd-380, 12'sd-1498, 12'sd-1200}},
{{12'sd-1325, 10'sd-368, 12'sd1035}, {12'sd-1958, 10'sd440, 10'sd336}, {11'sd579, 12'sd1304, 12'sd-1829}},
{{12'sd-1858, 11'sd517, 12'sd-1618}, {10'sd-428, 11'sd594, 12'sd1369}, {13'sd2512, 11'sd656, 12'sd1038}},
{{9'sd-166, 10'sd-391, 11'sd766}, {12'sd1644, 11'sd-884, 13'sd2492}, {11'sd-866, 9'sd137, 10'sd353}},
{{12'sd-1725, 13'sd2395, 9'sd-241}, {8'sd-112, 12'sd-1349, 12'sd-1419}, {12'sd1440, 13'sd2534, 10'sd-284}},
{{13'sd-2187, 13'sd2487, 12'sd-1358}, {9'sd-150, 13'sd3326, 11'sd-907}, {11'sd906, 12'sd1590, 13'sd-2772}}},
{
{{12'sd1738, 11'sd-668, 13'sd2452}, {11'sd-577, 12'sd1503, 12'sd-1453}, {12'sd-1403, 11'sd543, 11'sd-685}},
{{13'sd-2280, 13'sd2136, 11'sd521}, {12'sd-1903, 10'sd360, 9'sd-136}, {11'sd-642, 12'sd-1068, 11'sd-880}},
{{12'sd1920, 11'sd758, 13'sd2696}, {10'sd-357, 12'sd1756, 12'sd-1766}, {12'sd-1840, 12'sd-1688, 11'sd-599}},
{{13'sd3086, 13'sd-2080, 11'sd-787}, {11'sd1012, 12'sd1421, 10'sd312}, {12'sd1234, 11'sd-837, 11'sd-571}},
{{11'sd674, 11'sd-609, 5'sd-12}, {13'sd-2230, 12'sd-1956, 12'sd-1783}, {12'sd-1282, 13'sd-2345, 12'sd1192}},
{{9'sd202, 12'sd-1723, 5'sd10}, {9'sd183, 11'sd-909, 9'sd166}, {12'sd-1052, 8'sd74, 10'sd-293}},
{{12'sd-1370, 9'sd242, 13'sd3213}, {13'sd2301, 12'sd-1558, 12'sd-1685}, {13'sd2488, 10'sd-427, 12'sd1372}},
{{13'sd-2316, 10'sd-353, 13'sd-2298}, {9'sd-137, 13'sd3103, 11'sd-696}, {13'sd2470, 11'sd799, 11'sd-566}},
{{10'sd333, 13'sd2576, 12'sd-1736}, {13'sd-3421, 12'sd-1440, 11'sd768}, {12'sd-1543, 9'sd-252, 11'sd-826}},
{{13'sd-2758, 13'sd2131, 10'sd488}, {12'sd-1694, 11'sd-838, 10'sd503}, {10'sd496, 13'sd2558, 12'sd-1610}},
{{9'sd181, 7'sd-61, 12'sd1210}, {12'sd-1101, 12'sd-1970, 12'sd1731}, {13'sd2248, 12'sd-1411, 13'sd2692}},
{{13'sd-2511, 13'sd-2704, 10'sd-417}, {13'sd-2933, 12'sd-1143, 11'sd-702}, {12'sd1071, 4'sd5, 11'sd-992}},
{{11'sd-891, 12'sd1133, 11'sd800}, {13'sd-3107, 13'sd-3534, 13'sd2084}, {12'sd-1080, 12'sd1482, 10'sd-422}},
{{12'sd1654, 9'sd174, 13'sd-2918}, {13'sd2292, 12'sd-1552, 12'sd1263}, {12'sd1939, 8'sd-101, 12'sd-1182}},
{{11'sd-901, 12'sd1564, 11'sd-1000}, {9'sd-242, 13'sd2807, 10'sd-421}, {10'sd-438, 7'sd41, 11'sd-700}},
{{9'sd189, 12'sd-1682, 12'sd-1134}, {11'sd-768, 12'sd-1517, 12'sd1660}, {13'sd-2498, 11'sd805, 12'sd-1927}},
{{13'sd2379, 12'sd1056, 10'sd-423}, {13'sd-2382, 10'sd342, 12'sd1785}, {9'sd157, 12'sd1854, 12'sd1882}},
{{12'sd-1419, 12'sd1590, 12'sd-1338}, {11'sd-1017, 10'sd-465, 12'sd-1280}, {8'sd81, 13'sd-2961, 13'sd-4016}},
{{13'sd-2963, 13'sd-3079, 12'sd-1650}, {12'sd1241, 13'sd2499, 12'sd1364}, {13'sd-3091, 10'sd-317, 13'sd-3499}},
{{11'sd-891, 13'sd-2474, 10'sd475}, {12'sd1659, 9'sd206, 13'sd2530}, {13'sd2472, 13'sd2303, 11'sd728}},
{{14'sd4099, 12'sd1748, 13'sd2564}, {12'sd1714, 12'sd1668, 10'sd-393}, {10'sd411, 12'sd-1551, 13'sd2685}},
{{12'sd-1698, 13'sd-2904, 12'sd-1658}, {13'sd2085, 11'sd714, 9'sd199}, {12'sd-1301, 11'sd959, 11'sd-762}},
{{7'sd-57, 12'sd-1139, 11'sd618}, {10'sd257, 13'sd-2094, 10'sd-505}, {13'sd-2581, 11'sd-926, 10'sd434}},
{{11'sd597, 13'sd3122, 11'sd835}, {13'sd3142, 13'sd2742, 7'sd-57}, {10'sd-496, 10'sd-384, 11'sd786}},
{{12'sd-1767, 10'sd-494, 12'sd-1776}, {12'sd1285, 13'sd-2662, 10'sd472}, {10'sd400, 12'sd-1977, 11'sd-656}},
{{12'sd-1628, 11'sd-599, 13'sd2364}, {12'sd1509, 13'sd2432, 11'sd778}, {10'sd-290, 12'sd1062, 12'sd-1327}},
{{10'sd-403, 13'sd2101, 13'sd-2437}, {13'sd-2498, 11'sd-659, 11'sd846}, {13'sd2189, 13'sd2305, 11'sd683}},
{{14'sd-4458, 12'sd1339, 13'sd-2544}, {10'sd-332, 13'sd2315, 9'sd-139}, {12'sd1839, 13'sd-2496, 11'sd-943}},
{{12'sd-1126, 13'sd2420, 12'sd-1576}, {12'sd1089, 12'sd-1102, 12'sd-1965}, {11'sd-603, 10'sd-375, 12'sd-1296}},
{{11'sd787, 12'sd1734, 13'sd2980}, {11'sd-734, 9'sd195, 12'sd1464}, {11'sd965, 13'sd-2266, 11'sd589}},
{{13'sd3568, 12'sd-1938, 11'sd555}, {13'sd2528, 12'sd1492, 10'sd429}, {13'sd3933, 9'sd-172, 12'sd-1265}},
{{12'sd1067, 12'sd1818, 10'sd287}, {12'sd-1497, 13'sd-2283, 13'sd-2400}, {13'sd-2618, 13'sd2144, 11'sd-929}},
{{12'sd1387, 11'sd583, 13'sd-2329}, {11'sd704, 11'sd-945, 10'sd300}, {10'sd308, 11'sd-879, 11'sd518}},
{{11'sd-804, 12'sd1653, 9'sd131}, {10'sd-510, 12'sd1303, 12'sd-1372}, {13'sd-2064, 12'sd-1216, 12'sd1747}},
{{11'sd-887, 12'sd1157, 12'sd1543}, {11'sd-741, 11'sd-543, 13'sd-3080}, {12'sd-2025, 10'sd394, 13'sd-2112}},
{{11'sd-938, 11'sd-860, 13'sd2077}, {13'sd-3058, 12'sd-1395, 8'sd-92}, {11'sd670, 10'sd-298, 13'sd2081}},
{{13'sd-2168, 12'sd-1212, 12'sd1466}, {12'sd1463, 13'sd2894, 13'sd-2151}, {13'sd2209, 13'sd2966, 12'sd2018}},
{{11'sd-690, 10'sd-432, 12'sd1658}, {10'sd397, 12'sd-1226, 13'sd2242}, {12'sd1154, 13'sd2182, 12'sd1973}},
{{9'sd165, 12'sd1164, 12'sd1609}, {10'sd-346, 12'sd1527, 12'sd1077}, {12'sd1100, 5'sd-8, 11'sd847}},
{{12'sd-1137, 12'sd1532, 10'sd-283}, {11'sd-643, 13'sd-2167, 11'sd799}, {12'sd-1492, 13'sd2916, 10'sd-371}},
{{13'sd-3419, 10'sd-344, 12'sd-1769}, {10'sd369, 13'sd2192, 11'sd-845}, {11'sd778, 12'sd1715, 11'sd860}},
{{12'sd-1576, 11'sd676, 11'sd-935}, {12'sd-1297, 11'sd829, 11'sd-1002}, {12'sd1707, 11'sd-525, 13'sd2174}},
{{13'sd4004, 11'sd907, 12'sd1576}, {11'sd543, 11'sd574, 13'sd3057}, {10'sd348, 11'sd834, 12'sd1284}},
{{13'sd2765, 11'sd-733, 12'sd-1289}, {12'sd-1289, 12'sd-1692, 10'sd358}, {12'sd1379, 13'sd2410, 13'sd2382}},
{{8'sd-95, 12'sd1337, 12'sd-1499}, {13'sd3031, 11'sd-983, 12'sd-1254}, {8'sd117, 9'sd186, 10'sd-454}},
{{11'sd-1021, 13'sd2724, 8'sd109}, {9'sd-252, 12'sd-1817, 10'sd429}, {11'sd-983, 13'sd2452, 8'sd-76}},
{{13'sd2374, 12'sd1865, 13'sd2131}, {11'sd-757, 13'sd-2664, 13'sd-2485}, {10'sd-465, 10'sd470, 13'sd-2423}},
{{13'sd-2710, 12'sd-1359, 10'sd-500}, {9'sd-253, 13'sd-3085, 12'sd-1930}, {13'sd2417, 12'sd-1079, 12'sd1560}},
{{12'sd1435, 11'sd715, 12'sd-1214}, {13'sd3196, 13'sd2292, 10'sd-387}, {13'sd-2266, 12'sd1406, 11'sd928}},
{{12'sd-1430, 12'sd1984, 13'sd-3980}, {11'sd652, 11'sd-988, 10'sd-297}, {12'sd-1329, 9'sd225, 14'sd-4131}},
{{11'sd-779, 10'sd466, 11'sd-807}, {13'sd2183, 12'sd1124, 12'sd-1321}, {10'sd-375, 13'sd-2343, 13'sd-3209}},
{{12'sd1147, 12'sd-1763, 11'sd997}, {12'sd-1821, 12'sd-1864, 13'sd2228}, {12'sd1270, 12'sd1338, 13'sd2109}},
{{12'sd1087, 13'sd-2571, 11'sd-673}, {13'sd2868, 11'sd556, 12'sd-1747}, {11'sd1007, 11'sd-944, 12'sd1254}},
{{13'sd2757, 13'sd-2184, 13'sd-3325}, {11'sd538, 10'sd-342, 12'sd-1643}, {12'sd-1471, 10'sd-417, 12'sd-1168}},
{{13'sd3979, 10'sd433, 13'sd3679}, {13'sd2410, 11'sd-749, 10'sd355}, {12'sd1393, 13'sd-2303, 11'sd-871}},
{{12'sd-1653, 13'sd2787, 13'sd2630}, {12'sd1131, 11'sd-578, 12'sd1556}, {12'sd-1396, 11'sd850, 13'sd2395}},
{{11'sd742, 13'sd2132, 8'sd87}, {7'sd55, 12'sd1287, 13'sd2730}, {13'sd2850, 10'sd315, 12'sd-2046}},
{{10'sd-329, 13'sd2294, 12'sd-1593}, {13'sd-2133, 11'sd858, 13'sd-2869}, {12'sd1942, 12'sd1421, 10'sd-346}},
{{11'sd685, 13'sd-2856, 12'sd-1748}, {11'sd-696, 12'sd1186, 12'sd1075}, {13'sd3349, 12'sd2047, 12'sd-1178}},
{{13'sd2356, 10'sd-500, 9'sd241}, {12'sd-1422, 12'sd1070, 12'sd1329}, {12'sd1169, 13'sd2210, 13'sd2576}},
{{10'sd409, 12'sd1421, 12'sd-1209}, {10'sd473, 13'sd-2247, 13'sd-3213}, {12'sd1406, 13'sd2100, 12'sd1441}},
{{13'sd2114, 12'sd1751, 13'sd-2403}, {12'sd-1666, 12'sd-1995, 11'sd1006}, {13'sd3240, 10'sd295, 13'sd-3335}},
{{12'sd1580, 13'sd-3356, 9'sd-143}, {12'sd1285, 10'sd-453, 8'sd93}, {10'sd276, 12'sd-1838, 12'sd-1616}},
{{13'sd2926, 10'sd-264, 13'sd-2724}, {11'sd-994, 10'sd304, 11'sd-762}, {12'sd1487, 12'sd-1789, 12'sd-1628}}},
{
{{13'sd-3938, 13'sd-2103, 12'sd-1616}, {13'sd-3721, 13'sd-2429, 14'sd-4218}, {13'sd-3682, 12'sd1259, 11'sd-641}},
{{10'sd-266, 13'sd-2164, 13'sd-3190}, {11'sd-737, 12'sd-1417, 9'sd159}, {13'sd2282, 13'sd2299, 11'sd729}},
{{14'sd-5893, 11'sd-604, 12'sd-1581}, {14'sd-6286, 9'sd-157, 11'sd885}, {13'sd-2941, 12'sd1258, 10'sd-285}},
{{11'sd-724, 13'sd2216, 14'sd-4162}, {13'sd-3077, 11'sd-814, 11'sd783}, {11'sd619, 10'sd-294, 13'sd-3227}},
{{12'sd-1860, 11'sd-802, 10'sd-377}, {13'sd2329, 12'sd-1661, 13'sd2137}, {12'sd1024, 10'sd-288, 11'sd523}},
{{12'sd1878, 11'sd828, 12'sd1814}, {13'sd2150, 13'sd-2550, 9'sd-241}, {11'sd647, 11'sd-858, 11'sd696}},
{{12'sd-1757, 13'sd-2126, 13'sd2339}, {11'sd-983, 13'sd-3593, 12'sd-1861}, {13'sd-3918, 13'sd-3368, 13'sd-3625}},
{{13'sd-2784, 12'sd1850, 14'sd-5491}, {13'sd-2614, 10'sd495, 14'sd-5228}, {11'sd-684, 12'sd2026, 14'sd-4384}},
{{13'sd3870, 9'sd166, 11'sd817}, {12'sd1465, 11'sd-693, 9'sd195}, {8'sd87, 11'sd-609, 13'sd-2600}},
{{13'sd2056, 13'sd2553, 12'sd-1377}, {11'sd-794, 13'sd-2810, 12'sd-1040}, {13'sd-2150, 12'sd-1937, 7'sd46}},
{{11'sd777, 13'sd-2874, 13'sd2052}, {12'sd1060, 13'sd-2543, 11'sd-680}, {11'sd-643, 10'sd421, 12'sd1905}},
{{10'sd301, 13'sd-3013, 12'sd-1492}, {12'sd-1454, 12'sd-1139, 12'sd1575}, {12'sd-1388, 12'sd1974, 12'sd-1761}},
{{12'sd1201, 13'sd-2283, 12'sd1685}, {12'sd1692, 13'sd-3382, 7'sd-39}, {11'sd831, 11'sd-827, 11'sd519}},
{{13'sd-2678, 7'sd37, 11'sd589}, {13'sd2058, 13'sd-2274, 12'sd1183}, {11'sd527, 13'sd-2573, 11'sd839}},
{{13'sd3815, 10'sd317, 11'sd-572}, {12'sd2043, 11'sd-895, 13'sd2285}, {12'sd1358, 13'sd3646, 11'sd-929}},
{{12'sd1025, 12'sd-1076, 13'sd-3679}, {10'sd464, 8'sd73, 12'sd1570}, {12'sd-1504, 13'sd2153, 11'sd-970}},
{{12'sd-1041, 13'sd2076, 13'sd-3706}, {12'sd2003, 12'sd1524, 13'sd-2785}, {11'sd-788, 11'sd-877, 12'sd-1477}},
{{14'sd5522, 12'sd1501, 13'sd-2096}, {14'sd4206, 12'sd1686, 14'sd-4155}, {12'sd-1039, 5'sd-15, 12'sd-1256}},
{{11'sd697, 13'sd2075, 11'sd810}, {12'sd1737, 11'sd559, 11'sd631}, {10'sd366, 8'sd-103, 11'sd535}},
{{12'sd-1910, 11'sd-534, 11'sd-598}, {12'sd-1308, 13'sd-3065, 10'sd-271}, {12'sd-1267, 11'sd639, 13'sd-2215}},
{{13'sd-3063, 12'sd-1970, 13'sd-3208}, {13'sd-3886, 13'sd-2352, 11'sd-702}, {12'sd-1280, 13'sd-2532, 13'sd-4076}},
{{12'sd-1316, 13'sd-3552, 11'sd-905}, {9'sd132, 12'sd-1157, 11'sd590}, {10'sd376, 12'sd-1972, 13'sd2182}},
{{13'sd-2876, 12'sd1464, 13'sd-3364}, {12'sd-1239, 12'sd-1547, 13'sd-2799}, {11'sd-745, 12'sd-1209, 12'sd1044}},
{{12'sd1359, 12'sd1566, 12'sd1185}, {13'sd3377, 12'sd1365, 12'sd-1266}, {12'sd1284, 13'sd-2055, 12'sd-2017}},
{{11'sd719, 12'sd1246, 11'sd514}, {13'sd2088, 12'sd-1894, 13'sd2185}, {13'sd-3018, 11'sd-582, 11'sd-799}},
{{13'sd-2753, 12'sd1936, 11'sd923}, {11'sd-896, 12'sd-1364, 12'sd1217}, {11'sd-948, 12'sd-1566, 12'sd-1365}},
{{11'sd-977, 13'sd2420, 13'sd-2201}, {12'sd1761, 12'sd1333, 11'sd-792}, {12'sd-2029, 12'sd1371, 13'sd2545}},
{{11'sd802, 11'sd-628, 13'sd3034}, {14'sd4275, 12'sd-1423, 13'sd2933}, {13'sd2437, 13'sd-2953, 13'sd2512}},
{{13'sd-2806, 12'sd-1949, 14'sd5014}, {12'sd-1610, 12'sd1787, 14'sd5025}, {12'sd1590, 12'sd-1050, 11'sd560}},
{{12'sd-1869, 11'sd773, 8'sd-86}, {11'sd-525, 11'sd838, 13'sd-3419}, {11'sd991, 12'sd1860, 13'sd2685}},
{{12'sd1827, 10'sd-449, 12'sd1611}, {11'sd843, 13'sd2103, 12'sd-1839}, {14'sd4187, 8'sd-112, 11'sd1021}},
{{12'sd1052, 11'sd-658, 12'sd1381}, {10'sd-501, 8'sd-101, 10'sd-281}, {13'sd2354, 12'sd-1889, 7'sd-54}},
{{10'sd468, 12'sd-1158, 13'sd2669}, {13'sd-2191, 11'sd527, 10'sd475}, {10'sd-385, 13'sd2504, 12'sd1817}},
{{8'sd-109, 10'sd-435, 13'sd-3451}, {13'sd2378, 12'sd1317, 13'sd-3180}, {13'sd3590, 12'sd1269, 13'sd-2475}},
{{10'sd263, 11'sd913, 14'sd4346}, {13'sd-3942, 13'sd-2573, 12'sd-1153}, {13'sd-3152, 13'sd2165, 12'sd-1865}},
{{11'sd-873, 12'sd-1202, 12'sd1635}, {13'sd2590, 10'sd485, 13'sd2277}, {12'sd1382, 10'sd261, 12'sd1530}},
{{10'sd-294, 13'sd-2138, 13'sd2408}, {12'sd1044, 13'sd-3396, 13'sd-2583}, {12'sd1577, 13'sd-2538, 10'sd412}},
{{13'sd2283, 11'sd-525, 13'sd-2614}, {12'sd-1786, 13'sd-2761, 13'sd-2459}, {11'sd600, 10'sd465, 13'sd2271}},
{{11'sd752, 12'sd1561, 13'sd-3269}, {11'sd-985, 11'sd720, 8'sd-112}, {13'sd-2592, 12'sd1049, 11'sd749}},
{{13'sd2414, 13'sd-2318, 12'sd-1083}, {13'sd-2150, 13'sd2361, 12'sd-1757}, {11'sd-708, 12'sd-1168, 12'sd1028}},
{{13'sd2235, 12'sd-1056, 12'sd-1363}, {13'sd-3020, 13'sd-2352, 12'sd-1566}, {11'sd-755, 13'sd-2084, 13'sd2063}},
{{13'sd-2356, 11'sd792, 13'sd3552}, {12'sd-1180, 11'sd-883, 13'sd2332}, {10'sd-325, 13'sd-2423, 14'sd4403}},
{{12'sd-1264, 13'sd2147, 13'sd2585}, {13'sd-3418, 13'sd2199, 12'sd-1888}, {14'sd-5322, 13'sd-2626, 12'sd1976}},
{{12'sd-1781, 11'sd760, 11'sd574}, {12'sd1907, 8'sd76, 9'sd-157}, {10'sd-330, 9'sd-214, 11'sd-764}},
{{14'sd-6299, 12'sd-1955, 11'sd709}, {13'sd-4083, 12'sd1591, 13'sd2272}, {13'sd-3669, 12'sd-1338, 7'sd-48}},
{{12'sd1510, 12'sd1626, 13'sd-2429}, {9'sd174, 13'sd-2833, 12'sd-1639}, {13'sd-3095, 12'sd-1299, 12'sd1460}},
{{13'sd-2938, 12'sd1178, 13'sd2725}, {12'sd1269, 12'sd2047, 13'sd2702}, {11'sd-961, 13'sd-2768, 11'sd745}},
{{11'sd-640, 12'sd1956, 13'sd2918}, {13'sd-3759, 13'sd-2515, 11'sd950}, {13'sd2402, 11'sd897, 14'sd4640}},
{{14'sd4232, 12'sd-1973, 13'sd-2714}, {12'sd2013, 10'sd496, 14'sd-5135}, {11'sd906, 11'sd665, 13'sd-3442}},
{{14'sd7295, 12'sd1717, 13'sd2592}, {13'sd3913, 13'sd3858, 13'sd3635}, {14'sd4268, 10'sd334, 12'sd-1268}},
{{14'sd-4396, 11'sd-645, 10'sd268}, {13'sd-4069, 10'sd335, 14'sd5982}, {14'sd-6495, 13'sd-2300, 14'sd4274}},
{{13'sd-2795, 12'sd-1403, 12'sd1166}, {13'sd-2310, 11'sd829, 12'sd-1212}, {9'sd161, 13'sd-2543, 12'sd-1621}},
{{13'sd2965, 12'sd2031, 13'sd3522}, {10'sd402, 13'sd2819, 12'sd1994}, {12'sd1076, 13'sd2247, 11'sd584}},
{{11'sd-595, 11'sd-866, 11'sd-626}, {13'sd-2834, 13'sd2100, 8'sd96}, {13'sd-3130, 11'sd943, 13'sd-3596}},
{{13'sd-3300, 10'sd-350, 12'sd-1657}, {5'sd9, 10'sd470, 13'sd-3309}, {12'sd1263, 12'sd1601, 13'sd-2896}},
{{12'sd1193, 13'sd-2356, 11'sd868}, {4'sd-6, 10'sd-310, 12'sd1940}, {11'sd-764, 13'sd2239, 12'sd-1645}},
{{13'sd2140, 11'sd906, 7'sd44}, {13'sd-2688, 13'sd2120, 13'sd-2544}, {12'sd1346, 13'sd3469, 13'sd-2766}},
{{11'sd-960, 11'sd-733, 14'sd4309}, {11'sd696, 13'sd2056, 12'sd1811}, {12'sd-1753, 13'sd-2096, 13'sd-2188}},
{{12'sd-1139, 9'sd227, 12'sd1240}, {12'sd1816, 13'sd-2325, 11'sd-765}, {11'sd539, 12'sd1627, 12'sd-1159}},
{{13'sd-3827, 13'sd-2399, 8'sd83}, {8'sd94, 9'sd208, 10'sd-413}, {13'sd2707, 12'sd1695, 12'sd1410}},
{{9'sd-237, 9'sd-252, 13'sd-2328}, {13'sd3059, 10'sd340, 12'sd1209}, {11'sd631, 9'sd217, 13'sd2083}},
{{13'sd-3041, 13'sd2916, 13'sd-2089}, {12'sd-1204, 13'sd2155, 10'sd-380}, {14'sd-4479, 10'sd507, 9'sd248}},
{{13'sd-2216, 12'sd-1728, 12'sd1232}, {12'sd-1819, 13'sd2533, 9'sd-174}, {12'sd-1792, 8'sd115, 12'sd-1332}},
{{11'sd-744, 13'sd-3593, 12'sd-1769}, {11'sd-718, 9'sd-255, 12'sd-1389}, {12'sd-1734, 13'sd3424, 13'sd-2147}}},
{
{{9'sd-157, 12'sd-1156, 13'sd-2470}, {12'sd1402, 10'sd355, 12'sd-1161}, {13'sd-2108, 11'sd739, 13'sd2116}},
{{11'sd-806, 11'sd718, 12'sd1250}, {11'sd-708, 10'sd-300, 12'sd-2041}, {13'sd-2524, 11'sd949, 12'sd-1429}},
{{14'sd-4110, 13'sd-2321, 13'sd-4061}, {12'sd1238, 13'sd2803, 11'sd-845}, {10'sd-384, 11'sd654, 13'sd2491}},
{{11'sd-872, 13'sd-2279, 13'sd-2255}, {11'sd-534, 12'sd1971, 5'sd-9}, {8'sd-94, 12'sd-1059, 12'sd1319}},
{{12'sd-1634, 10'sd417, 12'sd1490}, {10'sd-280, 10'sd-501, 10'sd-456}, {12'sd-1648, 13'sd-2776, 11'sd670}},
{{13'sd2177, 12'sd-1364, 12'sd1732}, {8'sd-119, 12'sd1042, 12'sd1601}, {9'sd-129, 13'sd2188, 13'sd2483}},
{{12'sd2028, 13'sd2583, 12'sd1989}, {11'sd514, 11'sd891, 12'sd-1170}, {13'sd-2117, 11'sd-1011, 10'sd-314}},
{{10'sd362, 13'sd-2429, 12'sd1206}, {10'sd443, 10'sd-323, 13'sd-2893}, {11'sd601, 11'sd-737, 13'sd-2457}},
{{12'sd1624, 13'sd2158, 13'sd2896}, {12'sd-1141, 12'sd-1533, 9'sd222}, {12'sd1078, 13'sd2737, 13'sd3272}},
{{13'sd-2305, 10'sd285, 12'sd-1556}, {12'sd1946, 12'sd-1293, 5'sd-12}, {10'sd328, 12'sd1881, 11'sd-534}},
{{9'sd171, 13'sd2428, 12'sd-2028}, {12'sd-1629, 11'sd865, 12'sd-1193}, {12'sd1041, 13'sd2292, 12'sd1106}},
{{12'sd1996, 12'sd1505, 9'sd-246}, {12'sd1751, 11'sd-590, 9'sd246}, {12'sd1131, 12'sd1077, 13'sd2207}},
{{11'sd-907, 11'sd630, 12'sd1582}, {10'sd468, 13'sd2520, 13'sd2772}, {10'sd-308, 10'sd506, 12'sd1599}},
{{12'sd-2005, 12'sd1232, 12'sd-1215}, {12'sd-1157, 12'sd-1967, 11'sd-964}, {12'sd-1214, 13'sd-2482, 11'sd914}},
{{12'sd-1923, 12'sd-1084, 13'sd2290}, {13'sd2986, 13'sd2741, 12'sd1088}, {11'sd773, 12'sd1037, 12'sd1209}},
{{12'sd1030, 12'sd1096, 11'sd691}, {13'sd-2266, 11'sd579, 13'sd-2502}, {12'sd-1493, 10'sd-442, 12'sd-1442}},
{{13'sd-2326, 12'sd-1729, 12'sd-1226}, {13'sd-2509, 12'sd1746, 13'sd-2986}, {10'sd405, 9'sd-165, 13'sd-2855}},
{{12'sd-1844, 13'sd3111, 12'sd-1334}, {12'sd1696, 12'sd1939, 13'sd3011}, {11'sd-932, 13'sd-2062, 13'sd2179}},
{{11'sd-721, 13'sd2739, 12'sd-1723}, {12'sd-1417, 10'sd373, 12'sd-1293}, {9'sd-193, 12'sd-1099, 11'sd1009}},
{{11'sd531, 12'sd1988, 13'sd2776}, {11'sd-763, 12'sd1942, 12'sd-1791}, {13'sd-2323, 12'sd1245, 10'sd484}},
{{12'sd-1147, 12'sd1418, 13'sd2188}, {10'sd-354, 13'sd-2163, 11'sd897}, {12'sd-1473, 10'sd315, 13'sd-2050}},
{{12'sd1816, 11'sd-877, 13'sd-2600}, {12'sd-1341, 12'sd1066, 12'sd-1177}, {10'sd-322, 12'sd1507, 12'sd-1136}},
{{13'sd2072, 13'sd2257, 13'sd-2158}, {13'sd-2203, 11'sd717, 13'sd-2222}, {13'sd2561, 12'sd-1276, 12'sd-1431}},
{{7'sd32, 9'sd246, 12'sd1807}, {12'sd-1817, 11'sd-714, 12'sd1544}, {12'sd1612, 12'sd1450, 12'sd1818}},
{{12'sd-1459, 13'sd2657, 9'sd236}, {11'sd986, 13'sd2189, 10'sd-472}, {13'sd2368, 12'sd-1821, 12'sd1556}},
{{11'sd541, 12'sd1938, 13'sd-2407}, {12'sd2034, 12'sd1250, 12'sd1141}, {11'sd580, 12'sd-1408, 13'sd2251}},
{{5'sd-15, 12'sd1446, 13'sd2715}, {9'sd-138, 11'sd542, 12'sd1885}, {13'sd-2358, 12'sd1610, 13'sd2590}},
{{13'sd2786, 12'sd-1674, 7'sd-47}, {13'sd2529, 13'sd2574, 13'sd2767}, {11'sd981, 12'sd1574, 9'sd-234}},
{{13'sd-2290, 11'sd1022, 10'sd360}, {13'sd2630, 11'sd815, 11'sd565}, {12'sd1238, 13'sd2915, 12'sd1967}},
{{13'sd-2143, 13'sd-2237, 10'sd340}, {9'sd214, 11'sd-814, 13'sd-2248}, {12'sd1415, 11'sd-953, 13'sd2450}},
{{12'sd1671, 10'sd-307, 13'sd2310}, {12'sd-1106, 10'sd-467, 10'sd-456}, {11'sd-859, 12'sd-1435, 13'sd2268}},
{{11'sd938, 12'sd1917, 13'sd-2632}, {9'sd-233, 12'sd1985, 12'sd-1963}, {13'sd-2799, 12'sd-1732, 9'sd214}},
{{10'sd357, 13'sd-2093, 12'sd-1612}, {13'sd-2218, 12'sd2037, 10'sd411}, {11'sd987, 13'sd-2820, 13'sd2280}},
{{12'sd-1915, 12'sd1689, 12'sd-1354}, {12'sd1294, 12'sd1968, 13'sd-2048}, {12'sd-2036, 11'sd1009, 13'sd-3394}},
{{12'sd-1554, 13'sd2390, 12'sd1506}, {7'sd-42, 13'sd2667, 11'sd941}, {13'sd2466, 13'sd2787, 13'sd2328}},
{{11'sd722, 13'sd2919, 13'sd2779}, {11'sd982, 13'sd2675, 9'sd199}, {11'sd911, 12'sd-1742, 12'sd1479}},
{{10'sd499, 11'sd808, 12'sd1617}, {13'sd2058, 11'sd943, 10'sd-496}, {12'sd-1840, 13'sd-2324, 13'sd-2265}},
{{13'sd3017, 12'sd1447, 13'sd2736}, {12'sd1797, 12'sd-1255, 12'sd1426}, {11'sd-977, 12'sd-2014, 12'sd-1305}},
{{11'sd-753, 13'sd-3197, 9'sd245}, {11'sd539, 11'sd532, 8'sd87}, {13'sd2618, 12'sd1377, 11'sd735}},
{{12'sd-1040, 12'sd-1343, 4'sd-4}, {13'sd2221, 13'sd2175, 12'sd1973}, {11'sd634, 11'sd552, 11'sd-604}},
{{12'sd1458, 9'sd183, 13'sd2833}, {12'sd2008, 7'sd-59, 11'sd968}, {13'sd-2194, 9'sd145, 13'sd3044}},
{{11'sd-734, 13'sd-2080, 9'sd225}, {10'sd361, 12'sd1808, 12'sd1803}, {12'sd-1975, 10'sd447, 10'sd265}},
{{11'sd546, 12'sd-1560, 11'sd991}, {12'sd1961, 11'sd-955, 12'sd-1137}, {10'sd-376, 10'sd-419, 12'sd-1640}},
{{13'sd-2269, 13'sd-2214, 13'sd-2251}, {13'sd-2242, 12'sd-1223, 13'sd-2454}, {9'sd130, 7'sd50, 13'sd2257}},
{{11'sd555, 11'sd-882, 13'sd-2506}, {13'sd-2192, 11'sd-931, 10'sd-316}, {12'sd1787, 8'sd89, 5'sd15}},
{{9'sd-129, 10'sd-393, 12'sd-1106}, {8'sd67, 12'sd1294, 12'sd1662}, {12'sd1431, 13'sd2115, 9'sd-159}},
{{13'sd-2210, 9'sd204, 11'sd772}, {11'sd851, 13'sd3092, 12'sd-1837}, {11'sd-913, 13'sd2401, 12'sd1694}},
{{13'sd-2860, 13'sd-3168, 11'sd715}, {13'sd2291, 11'sd-541, 10'sd368}, {12'sd1635, 12'sd1706, 13'sd2746}},
{{11'sd1017, 8'sd92, 10'sd-483}, {9'sd-195, 13'sd-2789, 12'sd1080}, {13'sd-2530, 12'sd1115, 11'sd-626}},
{{12'sd1530, 9'sd-212, 12'sd-1355}, {11'sd-814, 12'sd2039, 11'sd-851}, {11'sd-648, 11'sd660, 12'sd1896}},
{{12'sd1601, 10'sd-506, 13'sd2629}, {13'sd-2785, 13'sd2266, 13'sd2261}, {13'sd-2189, 12'sd-1890, 12'sd-1277}},
{{13'sd-2556, 12'sd-1586, 12'sd-1693}, {10'sd-316, 9'sd158, 11'sd-1002}, {13'sd2229, 11'sd931, 12'sd-1087}},
{{12'sd1164, 9'sd-226, 13'sd-2284}, {12'sd-1114, 12'sd2034, 11'sd613}, {11'sd-747, 13'sd2440, 12'sd1495}},
{{13'sd2074, 12'sd1737, 12'sd1599}, {13'sd2140, 13'sd2544, 8'sd-90}, {13'sd-2063, 12'sd1321, 12'sd1749}},
{{9'sd-173, 13'sd-2252, 11'sd879}, {11'sd-888, 12'sd1434, 12'sd-1049}, {13'sd-2062, 13'sd2083, 12'sd1205}},
{{10'sd322, 12'sd1477, 13'sd2446}, {11'sd-755, 11'sd525, 13'sd2337}, {11'sd-852, 11'sd-717, 9'sd169}},
{{12'sd1559, 13'sd2371, 13'sd2229}, {12'sd1969, 10'sd-270, 12'sd-1550}, {11'sd749, 6'sd-21, 8'sd-66}},
{{12'sd-1531, 10'sd335, 12'sd-1538}, {13'sd2102, 12'sd-1469, 12'sd-1452}, {13'sd-2458, 13'sd2974, 12'sd1812}},
{{11'sd-739, 9'sd-232, 13'sd3108}, {13'sd2210, 7'sd45, 12'sd1112}, {9'sd168, 10'sd-464, 12'sd1996}},
{{12'sd-1834, 12'sd1513, 12'sd-1912}, {12'sd1280, 12'sd-1667, 11'sd606}, {11'sd658, 10'sd401, 12'sd2022}},
{{12'sd1198, 11'sd954, 12'sd-1366}, {12'sd1330, 13'sd-2827, 12'sd-1923}, {13'sd2090, 13'sd-2529, 10'sd-464}},
{{11'sd662, 8'sd-68, 12'sd-1053}, {12'sd-1820, 13'sd-2388, 13'sd-2260}, {12'sd1298, 13'sd-2535, 12'sd-1074}},
{{12'sd-1736, 12'sd-1090, 13'sd2297}, {12'sd-1513, 11'sd-965, 13'sd2087}, {12'sd1212, 13'sd2145, 11'sd-993}},
{{10'sd337, 13'sd-3087, 12'sd-2010}, {13'sd-2998, 10'sd-434, 10'sd-445}, {13'sd-2288, 12'sd1812, 11'sd832}}},
{
{{13'sd-2190, 11'sd-976, 11'sd783}, {12'sd1312, 13'sd-2248, 12'sd1706}, {12'sd1415, 11'sd987, 10'sd-317}},
{{12'sd-1526, 12'sd2032, 13'sd2346}, {11'sd-888, 10'sd-489, 11'sd-737}, {13'sd2136, 12'sd-2011, 10'sd-287}},
{{12'sd1144, 12'sd-1634, 10'sd-324}, {11'sd-1011, 10'sd-362, 11'sd999}, {12'sd1908, 13'sd3140, 11'sd-699}},
{{10'sd-351, 12'sd-1111, 10'sd498}, {13'sd2298, 8'sd102, 13'sd-2465}, {11'sd704, 11'sd807, 11'sd975}},
{{12'sd-1539, 11'sd874, 13'sd-2414}, {12'sd-1800, 11'sd828, 12'sd-1292}, {10'sd355, 10'sd364, 12'sd1542}},
{{11'sd903, 13'sd-2103, 11'sd796}, {12'sd-1195, 13'sd-2510, 11'sd558}, {12'sd1918, 13'sd2189, 13'sd2630}},
{{11'sd737, 12'sd1403, 12'sd-1288}, {11'sd880, 11'sd-769, 12'sd1391}, {12'sd1255, 13'sd-2568, 13'sd-2866}},
{{12'sd1793, 11'sd-592, 9'sd-208}, {11'sd-780, 13'sd2426, 8'sd-115}, {11'sd-791, 12'sd-1477, 11'sd835}},
{{12'sd-1047, 12'sd-1102, 12'sd-1341}, {9'sd-133, 13'sd2214, 11'sd-675}, {12'sd-1704, 12'sd-1935, 11'sd-647}},
{{13'sd2310, 11'sd1010, 12'sd1367}, {5'sd-10, 13'sd2626, 10'sd-362}, {7'sd54, 11'sd948, 12'sd1149}},
{{11'sd-971, 11'sd-519, 9'sd-213}, {12'sd1209, 11'sd705, 13'sd2685}, {13'sd-2555, 11'sd745, 11'sd-529}},
{{12'sd-1063, 12'sd1658, 12'sd1179}, {12'sd-1759, 9'sd219, 10'sd-469}, {12'sd1336, 13'sd-2141, 12'sd-1127}},
{{13'sd2485, 12'sd-1349, 9'sd-195}, {12'sd-1980, 11'sd579, 12'sd1323}, {12'sd-1402, 13'sd3797, 13'sd2259}},
{{13'sd-2077, 13'sd2545, 12'sd1554}, {12'sd1086, 12'sd-1996, 12'sd1181}, {12'sd-1235, 11'sd-913, 13'sd-2069}},
{{12'sd-1902, 11'sd686, 13'sd2477}, {11'sd786, 8'sd-81, 13'sd-2157}, {12'sd-1591, 11'sd-873, 13'sd-2107}},
{{12'sd1635, 13'sd2339, 10'sd291}, {10'sd-419, 12'sd-1525, 12'sd1662}, {13'sd3139, 11'sd560, 12'sd-1652}},
{{13'sd2150, 11'sd917, 13'sd-2547}, {13'sd-2467, 10'sd-472, 10'sd370}, {12'sd-1338, 11'sd955, 11'sd653}},
{{9'sd252, 13'sd-2300, 12'sd1683}, {7'sd37, 13'sd-2177, 11'sd-782}, {11'sd-916, 11'sd-698, 13'sd2242}},
{{11'sd-916, 13'sd-2328, 11'sd-863}, {12'sd1306, 13'sd-2288, 11'sd-676}, {12'sd-1502, 13'sd-2697, 12'sd-1032}},
{{11'sd923, 10'sd482, 10'sd-352}, {10'sd-486, 13'sd2691, 10'sd507}, {13'sd2271, 12'sd1381, 10'sd267}},
{{13'sd3323, 12'sd1173, 13'sd2903}, {12'sd1536, 12'sd1249, 12'sd1507}, {12'sd1518, 12'sd1152, 8'sd-92}},
{{13'sd-2739, 13'sd-2541, 13'sd2756}, {13'sd2597, 9'sd216, 12'sd-1922}, {11'sd-545, 12'sd1907, 12'sd-1627}},
{{12'sd1027, 12'sd1276, 12'sd1146}, {10'sd-436, 12'sd1074, 13'sd-2829}, {13'sd2571, 13'sd2163, 13'sd2236}},
{{13'sd2256, 11'sd-658, 13'sd-2385}, {12'sd-1863, 12'sd-1761, 12'sd2047}, {12'sd1580, 9'sd-225, 9'sd135}},
{{11'sd992, 13'sd2093, 12'sd2046}, {11'sd-836, 13'sd2937, 13'sd-2490}, {13'sd2479, 13'sd2515, 12'sd-1377}},
{{12'sd1112, 12'sd-1749, 12'sd-1314}, {12'sd1842, 10'sd-415, 8'sd-118}, {12'sd-1391, 7'sd45, 13'sd-2131}},
{{12'sd1412, 10'sd-409, 10'sd265}, {12'sd-1278, 11'sd563, 12'sd1572}, {12'sd-1906, 13'sd-2673, 11'sd-822}},
{{12'sd-1886, 12'sd1561, 11'sd-516}, {12'sd1250, 11'sd-591, 12'sd-1988}, {12'sd1761, 7'sd52, 13'sd-2596}},
{{11'sd-1020, 12'sd-1599, 13'sd-2216}, {12'sd1860, 13'sd2734, 13'sd2364}, {13'sd2947, 12'sd1615, 12'sd1638}},
{{11'sd-805, 8'sd78, 10'sd-293}, {13'sd-2453, 13'sd2322, 12'sd1908}, {12'sd1229, 12'sd-1052, 12'sd1375}},
{{11'sd-604, 10'sd472, 11'sd816}, {13'sd-2381, 9'sd-129, 8'sd71}, {12'sd1744, 11'sd-925, 13'sd-2699}},
{{12'sd1709, 8'sd-95, 11'sd769}, {12'sd-1119, 12'sd1477, 8'sd67}, {11'sd652, 12'sd1985, 13'sd-2521}},
{{10'sd-467, 12'sd-1714, 13'sd-3026}, {13'sd2576, 12'sd1686, 12'sd-1756}, {12'sd-1189, 11'sd-1004, 11'sd-675}},
{{13'sd2168, 12'sd1211, 13'sd-2083}, {12'sd-1836, 12'sd-1652, 12'sd-1191}, {13'sd-2697, 12'sd2005, 12'sd1157}},
{{13'sd2608, 12'sd1387, 9'sd-217}, {12'sd-1887, 9'sd184, 12'sd1146}, {12'sd-1081, 12'sd1260, 12'sd1326}},
{{12'sd-1185, 12'sd1457, 13'sd-2381}, {10'sd436, 9'sd-191, 12'sd1163}, {13'sd2599, 13'sd3009, 12'sd2045}},
{{12'sd-1298, 13'sd-2400, 11'sd620}, {11'sd-686, 12'sd1738, 13'sd2272}, {12'sd-1484, 12'sd-1532, 12'sd-1779}},
{{12'sd1740, 13'sd2456, 3'sd3}, {13'sd2492, 12'sd-1905, 11'sd-619}, {10'sd352, 12'sd1735, 13'sd-2125}},
{{12'sd1999, 10'sd-452, 12'sd-1643}, {13'sd-2428, 11'sd-814, 12'sd1255}, {12'sd1457, 13'sd-2278, 10'sd-503}},
{{12'sd-1038, 10'sd275, 11'sd534}, {10'sd319, 13'sd-2877, 12'sd2028}, {9'sd-230, 13'sd2208, 12'sd-1579}},
{{11'sd749, 13'sd3445, 12'sd1248}, {10'sd310, 10'sd509, 13'sd2589}, {12'sd-1543, 13'sd2904, 12'sd1967}},
{{11'sd-636, 13'sd-2189, 12'sd-1607}, {10'sd-267, 13'sd3151, 11'sd854}, {12'sd1337, 13'sd2386, 13'sd3311}},
{{13'sd3085, 13'sd-2076, 12'sd-1567}, {13'sd-2141, 12'sd1903, 11'sd-953}, {10'sd-344, 11'sd-952, 11'sd808}},
{{11'sd-607, 12'sd1654, 13'sd-2449}, {13'sd2857, 10'sd274, 12'sd1587}, {10'sd511, 12'sd1721, 11'sd-549}},
{{11'sd-684, 12'sd1697, 12'sd-1184}, {13'sd-2207, 12'sd1428, 12'sd1541}, {12'sd1182, 12'sd-1689, 12'sd-1848}},
{{13'sd-2621, 9'sd156, 12'sd-1456}, {11'sd-979, 13'sd2293, 13'sd-2172}, {13'sd2856, 12'sd1375, 13'sd-2183}},
{{11'sd-988, 12'sd-1866, 12'sd1919}, {10'sd483, 11'sd-805, 10'sd-306}, {12'sd-1251, 12'sd-1413, 11'sd516}},
{{9'sd184, 11'sd-1015, 13'sd3036}, {13'sd2598, 13'sd-2194, 11'sd941}, {10'sd441, 13'sd2864, 13'sd2049}},
{{9'sd188, 13'sd2949, 12'sd1961}, {13'sd-2666, 12'sd-1650, 12'sd1602}, {9'sd-187, 11'sd562, 11'sd-536}},
{{13'sd-2274, 12'sd1439, 9'sd172}, {12'sd-1508, 12'sd1444, 12'sd1234}, {12'sd1048, 11'sd-714, 13'sd-2780}},
{{11'sd-1007, 11'sd-521, 13'sd-2445}, {13'sd-2079, 12'sd1742, 10'sd359}, {13'sd-2572, 13'sd2075, 13'sd-3252}},
{{11'sd-572, 11'sd947, 12'sd1067}, {9'sd142, 10'sd493, 12'sd-1168}, {8'sd85, 11'sd-547, 12'sd1944}},
{{13'sd2222, 12'sd-1640, 11'sd-784}, {11'sd669, 9'sd136, 12'sd-1910}, {13'sd2364, 12'sd1555, 12'sd1027}},
{{12'sd-1279, 10'sd345, 10'sd396}, {11'sd637, 9'sd-241, 13'sd-2173}, {12'sd-1623, 12'sd-1411, 11'sd-977}},
{{9'sd-176, 11'sd761, 13'sd-2547}, {11'sd-627, 11'sd-621, 11'sd655}, {11'sd-805, 12'sd2018, 12'sd1520}},
{{9'sd140, 7'sd63, 12'sd1734}, {11'sd-630, 9'sd-210, 11'sd-903}, {11'sd875, 12'sd1506, 13'sd-2064}},
{{12'sd-1818, 12'sd1842, 10'sd435}, {12'sd-1639, 11'sd528, 11'sd-869}, {12'sd-1292, 13'sd-2177, 10'sd-375}},
{{9'sd206, 12'sd-1073, 13'sd2081}, {12'sd-1387, 9'sd238, 10'sd-364}, {12'sd1893, 13'sd-2624, 6'sd-30}},
{{11'sd-670, 12'sd1232, 11'sd-557}, {10'sd-394, 12'sd1732, 11'sd-584}, {10'sd-493, 12'sd1600, 10'sd484}},
{{11'sd624, 12'sd1344, 11'sd-660}, {11'sd809, 12'sd1398, 10'sd-418}, {12'sd1308, 10'sd-422, 13'sd3145}},
{{11'sd585, 11'sd725, 12'sd2026}, {7'sd-51, 12'sd-1547, 12'sd-1670}, {13'sd-2405, 12'sd2040, 12'sd-1250}},
{{11'sd-886, 13'sd2233, 13'sd-2302}, {11'sd-820, 13'sd2227, 13'sd-2442}, {9'sd189, 11'sd-942, 10'sd344}},
{{12'sd-1106, 13'sd-2081, 12'sd1088}, {13'sd-2174, 11'sd-707, 1'sd0}, {13'sd3369, 12'sd-1843, 12'sd1670}},
{{13'sd2132, 13'sd2151, 12'sd1686}, {12'sd-1868, 12'sd1285, 12'sd1909}, {11'sd-945, 8'sd124, 11'sd-606}}},
{
{{10'sd287, 11'sd-932, 10'sd434}, {11'sd-775, 11'sd869, 11'sd-876}, {13'sd-2884, 12'sd1806, 13'sd-2361}},
{{13'sd-2461, 13'sd-2318, 13'sd-2518}, {10'sd-470, 12'sd-1426, 12'sd-1098}, {13'sd2054, 13'sd-2833, 11'sd958}},
{{13'sd-2737, 9'sd-207, 12'sd-1897}, {13'sd2944, 11'sd800, 13'sd2362}, {12'sd-1868, 12'sd-1935, 13'sd-2434}},
{{12'sd1588, 12'sd1385, 11'sd1003}, {13'sd-2193, 10'sd-495, 9'sd147}, {13'sd-2326, 13'sd2545, 12'sd-1632}},
{{12'sd-1633, 12'sd1051, 12'sd1397}, {12'sd-1105, 12'sd-1059, 13'sd-2725}, {10'sd472, 13'sd2100, 13'sd2759}},
{{9'sd237, 12'sd2002, 12'sd1504}, {13'sd2740, 10'sd270, 12'sd1613}, {12'sd1231, 13'sd-2664, 9'sd-215}},
{{13'sd2754, 7'sd46, 12'sd1701}, {10'sd-338, 12'sd1070, 13'sd-2287}, {12'sd-1223, 13'sd-2798, 9'sd134}},
{{12'sd1605, 11'sd772, 12'sd-1438}, {11'sd-813, 13'sd-2210, 9'sd-155}, {11'sd-912, 10'sd-271, 12'sd1837}},
{{13'sd-2258, 13'sd-2269, 13'sd2297}, {11'sd-611, 9'sd214, 9'sd-215}, {13'sd3128, 11'sd-544, 13'sd2456}},
{{11'sd702, 13'sd2341, 10'sd410}, {7'sd60, 12'sd-1132, 12'sd-1931}, {12'sd1093, 12'sd1581, 12'sd1527}},
{{9'sd-190, 12'sd1740, 12'sd1849}, {12'sd1267, 10'sd-372, 13'sd3098}, {12'sd-1779, 12'sd-1368, 13'sd-2401}},
{{12'sd1549, 13'sd-2123, 10'sd-269}, {11'sd784, 12'sd-1107, 12'sd1871}, {12'sd-1917, 12'sd-1993, 11'sd771}},
{{13'sd3603, 11'sd533, 9'sd-149}, {13'sd2508, 11'sd-652, 12'sd1093}, {12'sd1168, 12'sd-1139, 13'sd-2290}},
{{11'sd795, 12'sd1275, 11'sd-995}, {11'sd672, 10'sd-434, 12'sd1107}, {13'sd-2701, 12'sd1739, 12'sd1515}},
{{12'sd1248, 12'sd-1656, 11'sd758}, {9'sd198, 7'sd60, 13'sd2249}, {13'sd2326, 13'sd2951, 11'sd900}},
{{11'sd683, 10'sd-380, 10'sd-379}, {13'sd-2581, 13'sd-2555, 11'sd683}, {10'sd323, 12'sd1781, 12'sd1502}},
{{13'sd2180, 12'sd-1671, 12'sd-1860}, {12'sd-1760, 12'sd1772, 12'sd1749}, {12'sd-1961, 10'sd326, 13'sd-2935}},
{{12'sd1107, 12'sd-1676, 10'sd-358}, {13'sd-2055, 13'sd2363, 13'sd2665}, {11'sd-531, 10'sd474, 12'sd1408}},
{{12'sd-1927, 13'sd2486, 12'sd1485}, {13'sd-2310, 9'sd-171, 12'sd1146}, {12'sd-1310, 8'sd-77, 12'sd1888}},
{{12'sd1922, 12'sd1818, 7'sd53}, {12'sd-1330, 11'sd852, 10'sd-465}, {13'sd2050, 13'sd2289, 10'sd271}},
{{13'sd-3466, 11'sd-1013, 11'sd648}, {12'sd1976, 10'sd437, 10'sd445}, {12'sd1057, 9'sd142, 12'sd-1469}},
{{12'sd1575, 13'sd2399, 12'sd1714}, {11'sd687, 13'sd2276, 13'sd2854}, {11'sd593, 11'sd-741, 12'sd-1677}},
{{12'sd-1219, 13'sd-2544, 11'sd996}, {8'sd98, 10'sd300, 13'sd-2068}, {13'sd-2107, 13'sd-2514, 11'sd595}},
{{10'sd-332, 9'sd217, 12'sd-1316}, {13'sd-3060, 6'sd19, 12'sd1760}, {13'sd-2746, 12'sd1288, 12'sd1299}},
{{10'sd385, 13'sd2570, 13'sd-2188}, {11'sd524, 13'sd2871, 12'sd1279}, {13'sd-2103, 13'sd2460, 11'sd667}},
{{9'sd174, 13'sd2983, 13'sd3021}, {13'sd-2256, 12'sd-1620, 11'sd600}, {10'sd-313, 9'sd-174, 12'sd1681}},
{{13'sd-2862, 13'sd-3011, 11'sd-835}, {13'sd-3148, 13'sd-2436, 13'sd-2393}, {13'sd2175, 12'sd1779, 13'sd-2145}},
{{11'sd-963, 12'sd1157, 12'sd-2025}, {13'sd-2539, 9'sd187, 12'sd-1466}, {13'sd-2854, 12'sd-1900, 12'sd-1398}},
{{10'sd-259, 11'sd875, 10'sd-473}, {13'sd-2381, 12'sd1904, 12'sd1098}, {8'sd-96, 12'sd-1208, 13'sd2368}},
{{11'sd763, 12'sd1787, 12'sd-1627}, {11'sd933, 8'sd76, 12'sd1419}, {13'sd-2225, 10'sd470, 11'sd722}},
{{12'sd1894, 12'sd1884, 13'sd2922}, {13'sd-3125, 13'sd3002, 9'sd245}, {11'sd-979, 12'sd-1489, 13'sd2114}},
{{13'sd-2989, 11'sd-757, 12'sd1246}, {12'sd1751, 8'sd99, 13'sd-2651}, {13'sd-2518, 12'sd-1390, 12'sd1618}},
{{12'sd1386, 12'sd-1181, 9'sd168}, {12'sd1209, 9'sd246, 10'sd307}, {11'sd-539, 13'sd2452, 13'sd2231}},
{{12'sd-1258, 9'sd211, 12'sd-1505}, {13'sd2473, 12'sd-1286, 12'sd1538}, {12'sd-1846, 11'sd868, 11'sd651}},
{{11'sd685, 13'sd2657, 12'sd-1195}, {12'sd-1842, 12'sd1397, 13'sd2802}, {13'sd2256, 11'sd818, 12'sd1676}},
{{11'sd-850, 12'sd-1126, 12'sd1070}, {10'sd457, 10'sd-509, 13'sd2811}, {11'sd-1000, 13'sd2847, 8'sd126}},
{{12'sd1435, 12'sd1878, 12'sd1444}, {12'sd1987, 13'sd2219, 12'sd1591}, {11'sd-647, 13'sd-2402, 13'sd-2342}},
{{13'sd2972, 12'sd1734, 13'sd2193}, {12'sd-1994, 8'sd-96, 13'sd2101}, {10'sd-358, 9'sd-220, 10'sd283}},
{{13'sd-2482, 11'sd1002, 11'sd-609}, {11'sd-590, 13'sd-2385, 13'sd-2900}, {13'sd2117, 13'sd-2188, 12'sd-1357}},
{{13'sd-2698, 12'sd-1489, 12'sd-2003}, {10'sd331, 12'sd1724, 10'sd-449}, {12'sd1951, 13'sd2086, 11'sd-650}},
{{12'sd1811, 11'sd790, 13'sd3019}, {12'sd1887, 12'sd1389, 13'sd2404}, {13'sd2729, 8'sd-76, 12'sd-1709}},
{{12'sd-1403, 10'sd480, 12'sd-1794}, {13'sd2329, 12'sd1891, 7'sd33}, {13'sd2635, 10'sd-319, 11'sd-725}},
{{12'sd1333, 10'sd405, 9'sd-211}, {9'sd243, 11'sd-726, 12'sd1383}, {11'sd-844, 13'sd-2112, 12'sd1149}},
{{12'sd1777, 13'sd3032, 12'sd1811}, {13'sd2910, 9'sd-182, 12'sd1371}, {11'sd525, 13'sd2234, 12'sd1331}},
{{12'sd-1533, 10'sd-397, 13'sd-2717}, {11'sd755, 12'sd1220, 12'sd1172}, {13'sd2511, 11'sd928, 12'sd1367}},
{{11'sd-950, 13'sd2685, 9'sd-139}, {13'sd-2121, 11'sd-836, 12'sd-1548}, {13'sd2567, 11'sd942, 12'sd1788}},
{{11'sd858, 13'sd2495, 10'sd-397}, {12'sd1716, 12'sd1245, 11'sd618}, {13'sd2354, 11'sd-978, 12'sd-1577}},
{{12'sd1282, 12'sd1956, 13'sd2772}, {6'sd31, 11'sd824, 13'sd-2500}, {10'sd504, 12'sd1540, 13'sd-2775}},
{{10'sd-502, 11'sd-977, 12'sd1316}, {9'sd-248, 12'sd1169, 12'sd-1595}, {10'sd-439, 12'sd-1200, 6'sd-24}},
{{10'sd-377, 9'sd-205, 12'sd1498}, {7'sd-45, 12'sd1251, 10'sd260}, {10'sd274, 13'sd2870, 13'sd2286}},
{{13'sd2221, 7'sd-32, 11'sd-792}, {13'sd-2297, 11'sd703, 12'sd-1943}, {13'sd2296, 12'sd-1478, 12'sd-1654}},
{{12'sd-1120, 13'sd2375, 12'sd-1638}, {12'sd-1578, 13'sd-2552, 10'sd325}, {12'sd1606, 13'sd2478, 11'sd-572}},
{{12'sd1478, 10'sd-511, 12'sd-1761}, {13'sd2306, 12'sd-1836, 12'sd-1460}, {12'sd1043, 13'sd2237, 12'sd-1805}},
{{9'sd140, 10'sd-509, 12'sd-1345}, {6'sd-16, 9'sd-193, 12'sd-1795}, {10'sd259, 9'sd-131, 13'sd2273}},
{{13'sd-2238, 12'sd1942, 12'sd-1786}, {13'sd-2087, 13'sd2906, 12'sd-1564}, {12'sd-1743, 10'sd-367, 12'sd2018}},
{{11'sd-777, 10'sd507, 13'sd2387}, {13'sd2991, 10'sd425, 11'sd-1011}, {11'sd-745, 13'sd-2418, 13'sd-2385}},
{{10'sd354, 11'sd-846, 12'sd-1282}, {13'sd-2278, 12'sd1768, 12'sd1794}, {11'sd-751, 9'sd-205, 13'sd-2415}},
{{12'sd-1780, 13'sd2650, 9'sd147}, {12'sd-1854, 11'sd-974, 12'sd-2031}, {8'sd-107, 9'sd-215, 13'sd2474}},
{{13'sd2499, 12'sd-1168, 9'sd-163}, {12'sd-1570, 12'sd1876, 12'sd1130}, {13'sd2073, 12'sd1793, 13'sd2481}},
{{11'sd651, 12'sd-1993, 13'sd-2503}, {11'sd-542, 11'sd714, 12'sd-1480}, {8'sd-115, 9'sd133, 12'sd-1418}},
{{12'sd-1292, 12'sd1781, 12'sd1909}, {13'sd-2808, 13'sd2053, 12'sd-1265}, {12'sd1399, 11'sd-801, 6'sd-25}},
{{8'sd91, 12'sd-1920, 12'sd1069}, {13'sd2254, 11'sd-945, 9'sd157}, {13'sd-2958, 12'sd1577, 12'sd-1745}},
{{8'sd97, 12'sd1094, 12'sd-1683}, {13'sd-2166, 11'sd-974, 10'sd-288}, {8'sd107, 13'sd2348, 11'sd682}},
{{13'sd-2860, 13'sd2429, 12'sd1859}, {13'sd-2306, 13'sd-2671, 12'sd-1073}, {12'sd1216, 11'sd965, 11'sd-558}}},
{
{{12'sd1186, 11'sd628, 11'sd811}, {10'sd-353, 12'sd-1289, 12'sd1756}, {12'sd1765, 9'sd-245, 12'sd1813}},
{{11'sd923, 13'sd-2131, 9'sd-253}, {13'sd2545, 13'sd-2452, 12'sd2042}, {11'sd-941, 11'sd630, 10'sd-381}},
{{7'sd-60, 11'sd611, 12'sd1961}, {12'sd1550, 8'sd-75, 4'sd5}, {13'sd-2334, 12'sd1788, 13'sd-2379}},
{{11'sd-518, 11'sd551, 7'sd-61}, {12'sd-1782, 12'sd-1761, 10'sd281}, {10'sd-432, 9'sd-179, 10'sd-266}},
{{12'sd-1131, 9'sd138, 12'sd2030}, {10'sd-491, 8'sd99, 12'sd1611}, {12'sd2025, 12'sd2040, 13'sd-2128}},
{{13'sd-2472, 12'sd1203, 13'sd-2824}, {9'sd-233, 11'sd-567, 13'sd-2160}, {6'sd29, 9'sd-178, 13'sd-2412}},
{{13'sd2293, 13'sd-2320, 12'sd-1411}, {13'sd2343, 12'sd1613, 10'sd316}, {11'sd-675, 13'sd-2935, 12'sd-2038}},
{{11'sd-585, 10'sd407, 7'sd-35}, {13'sd-2837, 11'sd880, 10'sd475}, {10'sd446, 13'sd2063, 12'sd1867}},
{{11'sd-580, 12'sd-1387, 12'sd-1611}, {9'sd155, 7'sd60, 13'sd-2731}, {8'sd79, 12'sd-1254, 12'sd1912}},
{{10'sd309, 12'sd1847, 11'sd701}, {13'sd-2050, 13'sd-2586, 12'sd-1442}, {12'sd1064, 13'sd-2128, 11'sd-540}},
{{13'sd2242, 8'sd-109, 11'sd662}, {12'sd1580, 9'sd-163, 13'sd2226}, {12'sd-1109, 11'sd818, 11'sd-670}},
{{12'sd1581, 11'sd-581, 10'sd-270}, {12'sd1327, 11'sd640, 12'sd1312}, {12'sd-1169, 12'sd-1810, 12'sd2035}},
{{12'sd1635, 11'sd883, 12'sd-1774}, {9'sd130, 13'sd-3528, 9'sd221}, {13'sd-3377, 13'sd-2350, 12'sd-1607}},
{{12'sd1367, 13'sd-2139, 13'sd2523}, {12'sd1281, 13'sd-2794, 11'sd819}, {12'sd-2003, 13'sd-2490, 12'sd1714}},
{{12'sd-1537, 13'sd-2611, 13'sd-2191}, {13'sd2622, 12'sd-2013, 13'sd2664}, {12'sd-1155, 11'sd-810, 13'sd2444}},
{{13'sd2529, 12'sd-1549, 12'sd-1265}, {13'sd-2206, 13'sd2571, 12'sd-1926}, {13'sd-2086, 12'sd-1756, 13'sd3225}},
{{12'sd-1567, 13'sd-2108, 12'sd-1798}, {11'sd-878, 10'sd-412, 12'sd1402}, {11'sd-658, 12'sd-1050, 12'sd1852}},
{{12'sd-1364, 12'sd1176, 9'sd216}, {13'sd-2132, 13'sd3772, 11'sd-827}, {13'sd-3281, 11'sd-985, 13'sd2623}},
{{12'sd1629, 10'sd-426, 12'sd1335}, {9'sd244, 12'sd-1703, 12'sd1321}, {10'sd275, 10'sd346, 12'sd-1196}},
{{10'sd-270, 12'sd-2004, 13'sd2816}, {13'sd-2271, 12'sd1107, 12'sd1686}, {13'sd2873, 9'sd172, 10'sd457}},
{{11'sd-981, 12'sd1437, 11'sd-957}, {11'sd822, 9'sd152, 12'sd1321}, {13'sd-2063, 12'sd1434, 12'sd1700}},
{{8'sd77, 13'sd-2852, 12'sd-1380}, {13'sd-2080, 10'sd370, 12'sd1489}, {10'sd419, 13'sd-2604, 12'sd1393}},
{{10'sd437, 12'sd1084, 8'sd96}, {11'sd701, 10'sd280, 12'sd-2019}, {11'sd624, 12'sd1410, 12'sd-1191}},
{{10'sd344, 12'sd-1515, 11'sd-549}, {10'sd375, 13'sd2599, 12'sd1288}, {13'sd-2861, 11'sd593, 12'sd1817}},
{{12'sd1253, 12'sd1278, 13'sd2684}, {12'sd1395, 12'sd-1743, 11'sd871}, {12'sd-1623, 13'sd-2252, 13'sd2468}},
{{12'sd1984, 11'sd-622, 12'sd1350}, {12'sd1805, 11'sd-618, 12'sd1064}, {13'sd-2055, 12'sd-2000, 12'sd1895}},
{{11'sd-908, 12'sd-1600, 13'sd-2389}, {13'sd-3048, 12'sd-1275, 13'sd-3160}, {12'sd1255, 11'sd572, 12'sd1836}},
{{8'sd-65, 12'sd1873, 11'sd-629}, {13'sd2376, 12'sd-1217, 13'sd-2051}, {10'sd387, 12'sd-1070, 11'sd-824}},
{{12'sd1325, 9'sd-255, 13'sd-2706}, {12'sd-1884, 9'sd189, 13'sd-2437}, {12'sd-1721, 10'sd-449, 11'sd711}},
{{11'sd568, 12'sd-1374, 11'sd768}, {13'sd-2119, 8'sd109, 13'sd-2648}, {9'sd241, 11'sd671, 10'sd479}},
{{10'sd-364, 14'sd4822, 8'sd-78}, {10'sd324, 13'sd2201, 11'sd697}, {11'sd553, 9'sd242, 11'sd955}},
{{13'sd-2673, 9'sd205, 11'sd-594}, {11'sd-639, 13'sd-2706, 10'sd-283}, {13'sd2496, 12'sd-1843, 12'sd-1663}},
{{11'sd-718, 11'sd-684, 11'sd872}, {11'sd925, 13'sd2729, 13'sd2511}, {13'sd-2628, 5'sd13, 13'sd2458}},
{{10'sd318, 11'sd-521, 11'sd931}, {12'sd1096, 11'sd949, 11'sd582}, {10'sd448, 13'sd-2058, 11'sd-595}},
{{12'sd1208, 12'sd1391, 11'sd-938}, {12'sd1543, 12'sd1597, 12'sd-1138}, {9'sd232, 11'sd-678, 13'sd-2182}},
{{11'sd-680, 12'sd-1481, 13'sd2674}, {11'sd-960, 13'sd2359, 10'sd459}, {12'sd1750, 11'sd545, 12'sd-1963}},
{{11'sd-577, 13'sd-2071, 9'sd-191}, {13'sd-2879, 10'sd356, 9'sd-209}, {12'sd1445, 11'sd-591, 6'sd-23}},
{{11'sd-818, 12'sd1602, 11'sd-567}, {13'sd2424, 12'sd1867, 13'sd-2261}, {12'sd1431, 11'sd-552, 13'sd2484}},
{{13'sd2211, 13'sd-2780, 12'sd1108}, {13'sd2480, 12'sd-1742, 12'sd1282}, {13'sd2660, 11'sd800, 12'sd1100}},
{{11'sd-1012, 11'sd-648, 12'sd1604}, {9'sd-228, 7'sd-52, 13'sd-2529}, {11'sd963, 12'sd1556, 12'sd-1320}},
{{11'sd629, 9'sd173, 12'sd1247}, {12'sd1678, 11'sd877, 12'sd1104}, {10'sd503, 12'sd-1188, 11'sd755}},
{{12'sd1810, 11'sd-537, 12'sd1916}, {13'sd2219, 12'sd-1284, 10'sd414}, {13'sd-2389, 12'sd-1536, 10'sd-333}},
{{11'sd-590, 13'sd-2115, 13'sd-2335}, {12'sd1684, 11'sd-617, 13'sd-2495}, {13'sd-2375, 12'sd1600, 13'sd-2238}},
{{12'sd-2026, 12'sd-1617, 12'sd1560}, {8'sd-100, 12'sd-1467, 12'sd-1607}, {11'sd916, 13'sd2802, 12'sd1038}},
{{13'sd-2245, 12'sd1027, 13'sd-2636}, {13'sd2693, 12'sd1668, 12'sd1221}, {9'sd-235, 12'sd-1137, 10'sd341}},
{{12'sd1710, 11'sd-780, 11'sd-775}, {7'sd-62, 11'sd564, 12'sd2036}, {11'sd671, 13'sd2852, 13'sd2366}},
{{12'sd1871, 12'sd1469, 13'sd2689}, {13'sd-2154, 13'sd2948, 11'sd870}, {10'sd-410, 11'sd-707, 5'sd-11}},
{{11'sd595, 13'sd-2190, 8'sd70}, {13'sd2488, 12'sd-1854, 12'sd1297}, {13'sd-2292, 13'sd-3494, 9'sd228}},
{{13'sd-3714, 13'sd2236, 13'sd2996}, {12'sd1362, 11'sd-751, 12'sd-1234}, {12'sd-2038, 13'sd2861, 8'sd96}},
{{13'sd-2958, 9'sd147, 11'sd852}, {12'sd-1537, 12'sd1294, 5'sd11}, {13'sd-3192, 13'sd3398, 13'sd2619}},
{{13'sd3175, 12'sd-1223, 12'sd1482}, {13'sd3694, 12'sd-1564, 11'sd591}, {11'sd649, 11'sd-728, 8'sd100}},
{{9'sd-215, 12'sd1109, 11'sd-875}, {12'sd1831, 11'sd-979, 12'sd-1754}, {11'sd698, 11'sd-837, 12'sd-1446}},
{{11'sd-655, 11'sd913, 13'sd2552}, {10'sd-270, 11'sd-797, 11'sd642}, {12'sd1170, 11'sd-818, 13'sd2353}},
{{12'sd1617, 10'sd302, 12'sd1119}, {13'sd-2372, 12'sd1825, 13'sd-2390}, {10'sd-343, 10'sd427, 6'sd22}},
{{13'sd3216, 12'sd1188, 12'sd1541}, {11'sd940, 9'sd-252, 12'sd1053}, {10'sd-458, 13'sd-2075, 11'sd932}},
{{13'sd-2484, 11'sd-946, 13'sd2767}, {12'sd1721, 9'sd-217, 11'sd878}, {10'sd312, 9'sd-165, 13'sd-2727}},
{{9'sd-200, 12'sd1966, 13'sd2255}, {13'sd-2271, 13'sd2770, 11'sd-951}, {11'sd-619, 12'sd-1559, 11'sd-774}},
{{11'sd-814, 12'sd-1750, 13'sd2417}, {11'sd540, 11'sd583, 10'sd-417}, {13'sd-2849, 11'sd-791, 11'sd612}},
{{8'sd-126, 12'sd1135, 13'sd3277}, {12'sd1712, 11'sd528, 12'sd1513}, {13'sd-2455, 13'sd-2351, 12'sd1077}},
{{12'sd-1912, 13'sd2373, 12'sd-1949}, {11'sd-602, 10'sd-326, 12'sd-1822}, {13'sd-2838, 9'sd211, 13'sd-2913}},
{{10'sd-310, 8'sd-120, 11'sd-969}, {10'sd-352, 11'sd-648, 12'sd-1839}, {13'sd-2200, 8'sd125, 11'sd860}},
{{8'sd94, 12'sd-1575, 12'sd1513}, {11'sd-591, 12'sd1569, 12'sd-1424}, {12'sd1957, 13'sd-2471, 12'sd1213}},
{{13'sd-2129, 11'sd908, 12'sd1102}, {12'sd-1630, 12'sd-1153, 12'sd-1187}, {9'sd213, 13'sd2558, 12'sd1095}},
{{13'sd-2317, 11'sd-742, 13'sd2492}, {13'sd2726, 12'sd-1784, 7'sd37}, {11'sd-891, 13'sd2408, 8'sd-91}}},
{
{{12'sd1747, 12'sd1383, 11'sd964}, {12'sd1468, 13'sd2199, 13'sd2950}, {12'sd2016, 12'sd-1308, 9'sd-154}},
{{12'sd1613, 12'sd-2005, 11'sd722}, {13'sd-2945, 12'sd-1511, 11'sd-864}, {12'sd-1789, 8'sd-105, 11'sd979}},
{{14'sd4921, 11'sd891, 13'sd2623}, {13'sd-2342, 9'sd187, 11'sd972}, {12'sd-1211, 11'sd992, 10'sd455}},
{{12'sd-1469, 13'sd-2514, 13'sd-2743}, {11'sd728, 11'sd-985, 8'sd74}, {12'sd-1815, 12'sd1302, 12'sd-1705}},
{{11'sd542, 13'sd2090, 8'sd78}, {12'sd-1119, 12'sd1549, 13'sd2321}, {11'sd737, 10'sd-372, 13'sd2514}},
{{11'sd-861, 10'sd420, 12'sd-1944}, {13'sd2175, 12'sd-1996, 9'sd-132}, {11'sd559, 11'sd867, 12'sd2034}},
{{12'sd-1162, 13'sd2397, 11'sd-1010}, {13'sd2300, 12'sd-1760, 9'sd148}, {9'sd-156, 13'sd2490, 13'sd-2887}},
{{10'sd401, 12'sd-1844, 11'sd-780}, {13'sd-2654, 11'sd-939, 12'sd-1466}, {11'sd805, 12'sd-1155, 13'sd-2615}},
{{13'sd2573, 13'sd-2336, 13'sd2611}, {10'sd280, 10'sd301, 11'sd-1010}, {14'sd4776, 10'sd-466, 12'sd-1405}},
{{12'sd-1930, 13'sd2440, 13'sd-2067}, {12'sd-2015, 12'sd1412, 12'sd-1497}, {12'sd-1044, 13'sd-2448, 12'sd-1549}},
{{13'sd-2157, 9'sd240, 13'sd2324}, {12'sd1332, 9'sd206, 10'sd342}, {11'sd903, 12'sd-1168, 10'sd-495}},
{{11'sd-969, 8'sd64, 12'sd-1107}, {3'sd2, 12'sd-1945, 12'sd1645}, {13'sd-2168, 12'sd-1332, 12'sd1585}},
{{8'sd-94, 13'sd2361, 11'sd633}, {8'sd120, 11'sd-929, 10'sd340}, {8'sd-111, 8'sd-87, 10'sd-372}},
{{12'sd-1373, 11'sd-700, 12'sd-1964}, {12'sd-1533, 12'sd-1769, 12'sd-1855}, {13'sd-2933, 11'sd-655, 12'sd1177}},
{{11'sd681, 13'sd-2731, 10'sd-303}, {10'sd416, 13'sd2887, 10'sd339}, {9'sd177, 12'sd-1060, 12'sd1415}},
{{12'sd-1214, 12'sd-1339, 12'sd-2022}, {12'sd-1581, 13'sd2163, 13'sd2479}, {12'sd-1600, 10'sd-417, 11'sd633}},
{{12'sd2021, 12'sd-1681, 12'sd-1634}, {12'sd1769, 12'sd1949, 12'sd1538}, {12'sd1933, 10'sd393, 11'sd736}},
{{12'sd1179, 12'sd-1306, 13'sd-3260}, {9'sd-182, 11'sd-532, 12'sd-2016}, {12'sd-1822, 13'sd-2461, 13'sd2425}},
{{9'sd-169, 10'sd-461, 11'sd-977}, {13'sd2398, 12'sd-1176, 13'sd3076}, {12'sd-1862, 13'sd-3168, 9'sd-170}},
{{7'sd48, 12'sd1790, 11'sd743}, {12'sd-1348, 10'sd-267, 13'sd2208}, {11'sd-959, 11'sd-926, 11'sd-774}},
{{11'sd669, 13'sd2061, 13'sd2067}, {13'sd-2604, 13'sd-2091, 13'sd-2410}, {14'sd4974, 13'sd3264, 12'sd1105}},
{{10'sd314, 10'sd-285, 11'sd-853}, {12'sd-1100, 12'sd1101, 12'sd-1033}, {12'sd1899, 13'sd-2626, 10'sd391}},
{{10'sd328, 12'sd-1447, 12'sd1618}, {11'sd609, 13'sd2456, 13'sd-2727}, {12'sd1654, 13'sd2058, 9'sd-240}},
{{10'sd314, 12'sd1594, 11'sd583}, {8'sd-126, 12'sd-1058, 13'sd-2511}, {8'sd-66, 12'sd1702, 13'sd2338}},
{{12'sd-1600, 13'sd-2868, 12'sd-1221}, {11'sd919, 12'sd1884, 13'sd2912}, {12'sd-2035, 13'sd-2436, 13'sd-2346}},
{{6'sd-19, 11'sd623, 12'sd-1703}, {12'sd-1779, 13'sd-2502, 12'sd1548}, {13'sd2829, 12'sd-2044, 9'sd165}},
{{11'sd-686, 13'sd2215, 12'sd1285}, {13'sd-2305, 12'sd1713, 10'sd-256}, {13'sd-2640, 12'sd-1803, 13'sd2118}},
{{13'sd-2933, 13'sd-2359, 13'sd3072}, {12'sd1987, 13'sd-2086, 11'sd-990}, {5'sd-10, 11'sd-860, 10'sd-413}},
{{8'sd76, 12'sd-2028, 13'sd2978}, {11'sd-808, 12'sd-1399, 12'sd1304}, {12'sd1820, 10'sd294, 12'sd1894}},
{{8'sd124, 8'sd66, 13'sd-3276}, {10'sd-275, 13'sd-2246, 12'sd-1571}, {11'sd650, 10'sd-259, 12'sd1524}},
{{12'sd1395, 11'sd728, 10'sd369}, {13'sd-2403, 13'sd-3663, 7'sd46}, {12'sd-1784, 13'sd-2837, 13'sd-3457}},
{{11'sd855, 13'sd3188, 11'sd605}, {11'sd586, 13'sd-2259, 13'sd2301}, {12'sd1339, 13'sd2642, 10'sd-471}},
{{13'sd-2247, 9'sd150, 12'sd1799}, {13'sd-2791, 11'sd670, 9'sd254}, {10'sd-396, 10'sd-482, 12'sd1063}},
{{10'sd390, 13'sd2641, 12'sd1981}, {12'sd-2012, 11'sd987, 13'sd-2478}, {11'sd621, 10'sd-490, 6'sd19}},
{{9'sd-142, 10'sd-397, 11'sd775}, {11'sd836, 12'sd-1168, 11'sd-534}, {7'sd61, 12'sd2002, 12'sd-1194}},
{{13'sd-2734, 12'sd-1136, 13'sd-2146}, {13'sd2552, 12'sd1891, 13'sd-2820}, {13'sd2499, 10'sd-368, 11'sd-770}},
{{12'sd-1985, 6'sd-20, 12'sd1302}, {12'sd-1060, 12'sd-1151, 13'sd-2696}, {12'sd-1505, 13'sd-2398, 9'sd128}},
{{8'sd89, 12'sd1600, 11'sd-686}, {12'sd1435, 12'sd1551, 11'sd811}, {10'sd375, 11'sd-971, 12'sd1947}},
{{12'sd2022, 10'sd-371, 8'sd-125}, {11'sd953, 12'sd1371, 13'sd2291}, {12'sd-1571, 10'sd443, 12'sd1809}},
{{11'sd-686, 13'sd-2163, 12'sd-1815}, {12'sd1772, 8'sd65, 9'sd-148}, {13'sd-2292, 10'sd350, 13'sd-3113}},
{{7'sd-51, 11'sd-926, 11'sd-766}, {13'sd3075, 11'sd-911, 13'sd-2440}, {13'sd2584, 10'sd500, 12'sd-1476}},
{{12'sd-1220, 11'sd544, 8'sd-101}, {13'sd-3591, 11'sd-1005, 12'sd1885}, {13'sd-2794, 12'sd1824, 12'sd1461}},
{{10'sd397, 8'sd-80, 13'sd2711}, {12'sd-1825, 11'sd-806, 12'sd-1598}, {13'sd2438, 12'sd1228, 13'sd3739}},
{{12'sd1405, 12'sd1217, 10'sd410}, {12'sd2021, 12'sd1235, 9'sd-147}, {12'sd1675, 13'sd2124, 11'sd833}},
{{14'sd4696, 11'sd987, 10'sd-329}, {11'sd754, 9'sd162, 11'sd846}, {12'sd1498, 12'sd1710, 13'sd-2088}},
{{11'sd-704, 8'sd78, 6'sd29}, {12'sd1658, 12'sd-1351, 7'sd35}, {13'sd2776, 13'sd2826, 12'sd1072}},
{{13'sd2095, 13'sd-2079, 11'sd-775}, {12'sd-1938, 13'sd-2554, 10'sd-455}, {11'sd766, 11'sd832, 11'sd897}},
{{14'sd4824, 10'sd475, 12'sd1795}, {12'sd-1050, 12'sd-1483, 10'sd412}, {13'sd-2155, 12'sd-1614, 12'sd-1722}},
{{12'sd1066, 13'sd2056, 9'sd-251}, {12'sd1860, 12'sd1216, 13'sd-2333}, {12'sd1432, 12'sd-1081, 12'sd-1984}},
{{12'sd-1500, 13'sd-3257, 9'sd244}, {13'sd2934, 12'sd1817, 13'sd3717}, {12'sd-1524, 12'sd-1345, 12'sd-1675}},
{{10'sd-269, 10'sd-457, 9'sd166}, {11'sd-752, 12'sd1602, 10'sd-272}, {13'sd2576, 13'sd-2179, 7'sd-63}},
{{11'sd637, 13'sd2888, 8'sd-68}, {9'sd-246, 12'sd-1507, 11'sd836}, {13'sd-2118, 11'sd-835, 9'sd210}},
{{10'sd-357, 13'sd-2616, 11'sd907}, {10'sd504, 13'sd-3099, 12'sd1046}, {12'sd1413, 11'sd-1006, 6'sd17}},
{{9'sd221, 10'sd-469, 12'sd1562}, {11'sd844, 12'sd-1638, 12'sd-1889}, {8'sd-80, 10'sd-511, 12'sd-1528}},
{{13'sd-2168, 12'sd1703, 9'sd217}, {11'sd-794, 12'sd-1280, 11'sd606}, {12'sd-1668, 10'sd-335, 13'sd2761}},
{{13'sd3429, 13'sd-2054, 12'sd-1769}, {12'sd1341, 11'sd528, 12'sd-1589}, {13'sd2161, 12'sd1949, 12'sd-1262}},
{{12'sd1567, 13'sd2823, 12'sd-1178}, {8'sd65, 11'sd-633, 7'sd34}, {12'sd1039, 13'sd-3085, 11'sd-1018}},
{{12'sd-1279, 11'sd644, 11'sd-573}, {13'sd-2227, 13'sd2233, 10'sd-476}, {8'sd117, 13'sd2173, 10'sd293}},
{{12'sd-1379, 11'sd-648, 13'sd-2056}, {13'sd-2606, 8'sd113, 13'sd-2447}, {12'sd-1260, 13'sd2088, 10'sd379}},
{{12'sd-1112, 10'sd280, 13'sd3870}, {12'sd-1042, 8'sd126, 12'sd1567}, {12'sd1432, 13'sd-2179, 11'sd-655}},
{{11'sd1003, 8'sd65, 11'sd882}, {12'sd-1190, 12'sd1641, 11'sd639}, {13'sd2167, 11'sd590, 13'sd-2978}},
{{13'sd-2827, 13'sd-2355, 9'sd-151}, {11'sd-741, 11'sd-952, 12'sd-1663}, {12'sd1227, 12'sd1932, 13'sd-2787}},
{{12'sd-2009, 13'sd-2066, 11'sd-855}, {7'sd-42, 12'sd1681, 12'sd1956}, {13'sd-4066, 11'sd525, 11'sd651}},
{{12'sd1300, 12'sd-1789, 12'sd1307}, {11'sd702, 9'sd-209, 11'sd-798}, {13'sd2050, 6'sd16, 13'sd-3182}}},
{
{{13'sd-2802, 11'sd744, 10'sd-408}, {12'sd-1714, 13'sd-2987, 13'sd2979}, {9'sd-227, 11'sd-950, 12'sd1716}},
{{11'sd854, 12'sd-1062, 12'sd1060}, {13'sd2222, 12'sd1567, 10'sd-319}, {11'sd-801, 9'sd156, 13'sd-2216}},
{{13'sd-3174, 12'sd-1028, 9'sd-253}, {13'sd-3005, 13'sd-3522, 11'sd1017}, {11'sd714, 12'sd-1163, 12'sd1296}},
{{13'sd3208, 11'sd-660, 13'sd3344}, {12'sd-1753, 12'sd-1531, 6'sd-19}, {13'sd2204, 12'sd-1845, 13'sd3341}},
{{13'sd-2484, 11'sd1011, 12'sd1770}, {12'sd1971, 12'sd1504, 12'sd-1625}, {11'sd-889, 10'sd-303, 13'sd2382}},
{{13'sd2680, 12'sd-1726, 13'sd-3084}, {7'sd51, 7'sd-59, 12'sd1583}, {5'sd-10, 12'sd1104, 12'sd1131}},
{{12'sd1620, 13'sd2673, 11'sd-666}, {13'sd-2446, 12'sd1556, 13'sd-2849}, {13'sd-2554, 12'sd1190, 12'sd-1715}},
{{10'sd-484, 13'sd-2500, 8'sd112}, {9'sd-243, 12'sd1819, 10'sd-319}, {6'sd25, 12'sd-1633, 11'sd-719}},
{{11'sd737, 13'sd-2072, 11'sd-645}, {12'sd1977, 13'sd-2068, 13'sd2314}, {12'sd1792, 12'sd-1634, 11'sd-565}},
{{12'sd-1952, 10'sd-434, 11'sd-552}, {13'sd-2350, 12'sd-1167, 13'sd-3336}, {12'sd-1923, 10'sd463, 11'sd797}},
{{13'sd-2616, 11'sd976, 9'sd-219}, {11'sd-880, 12'sd-1397, 10'sd331}, {12'sd-1392, 13'sd2541, 12'sd1667}},
{{12'sd-1087, 11'sd-900, 12'sd1348}, {12'sd1185, 12'sd1389, 12'sd-1850}, {13'sd-2900, 8'sd-76, 13'sd-2349}},
{{11'sd-801, 13'sd-2677, 12'sd1122}, {13'sd2921, 8'sd117, 9'sd204}, {11'sd826, 7'sd-59, 9'sd-130}},
{{8'sd118, 12'sd-1147, 11'sd-542}, {12'sd1928, 13'sd-2720, 12'sd-1881}, {13'sd-2537, 9'sd-252, 11'sd-565}},
{{12'sd1286, 13'sd3075, 12'sd1308}, {13'sd2696, 13'sd-2323, 11'sd782}, {13'sd3355, 8'sd90, 13'sd2883}},
{{11'sd-648, 13'sd2945, 12'sd1562}, {12'sd-1950, 12'sd1995, 11'sd-520}, {11'sd-757, 12'sd1304, 11'sd-805}},
{{12'sd1063, 10'sd-465, 10'sd-369}, {10'sd434, 12'sd1855, 12'sd-1764}, {10'sd-400, 13'sd2182, 12'sd1109}},
{{11'sd543, 12'sd-1474, 12'sd-1083}, {11'sd700, 12'sd-1575, 13'sd3365}, {10'sd-464, 13'sd-2344, 13'sd2447}},
{{12'sd1889, 13'sd3511, 12'sd1045}, {11'sd893, 13'sd-2050, 13'sd2397}, {12'sd-1654, 11'sd-981, 8'sd-108}},
{{12'sd-1351, 11'sd734, 11'sd567}, {12'sd-1540, 12'sd1641, 11'sd-915}, {11'sd689, 13'sd-2299, 8'sd93}},
{{12'sd-1915, 10'sd301, 13'sd-3841}, {13'sd-3308, 9'sd-162, 9'sd-233}, {14'sd-5922, 13'sd-2809, 11'sd-848}},
{{11'sd651, 12'sd-1359, 12'sd-1175}, {13'sd2766, 7'sd62, 9'sd-222}, {12'sd1544, 12'sd1547, 11'sd771}},
{{11'sd707, 12'sd-1710, 12'sd-1487}, {10'sd307, 10'sd-496, 11'sd-732}, {12'sd-1095, 11'sd541, 12'sd1321}},
{{13'sd-2132, 12'sd-1791, 12'sd1794}, {13'sd3337, 11'sd-726, 11'sd-678}, {13'sd3173, 12'sd-1750, 12'sd1695}},
{{11'sd1011, 10'sd317, 12'sd1896}, {9'sd-182, 12'sd1059, 12'sd1351}, {10'sd367, 12'sd-1244, 12'sd-1431}},
{{12'sd-1592, 13'sd2059, 12'sd1946}, {11'sd721, 13'sd2780, 12'sd1155}, {13'sd2588, 12'sd1849, 9'sd156}},
{{13'sd2432, 12'sd1442, 10'sd349}, {11'sd652, 12'sd-1367, 9'sd-210}, {12'sd1356, 13'sd2816, 10'sd363}},
{{13'sd2192, 10'sd313, 12'sd-1652}, {10'sd356, 11'sd592, 13'sd2289}, {10'sd-411, 13'sd2394, 7'sd-59}},
{{12'sd-1724, 13'sd2777, 12'sd1046}, {9'sd-135, 13'sd-2512, 12'sd1833}, {13'sd2885, 12'sd-1790, 12'sd1905}},
{{12'sd-1366, 12'sd1560, 13'sd2171}, {13'sd2150, 12'sd1075, 11'sd-608}, {11'sd-925, 11'sd-867, 12'sd-1951}},
{{11'sd-590, 10'sd-489, 10'sd-322}, {12'sd-1494, 13'sd-2421, 10'sd310}, {10'sd316, 11'sd675, 12'sd-1034}},
{{13'sd-3221, 10'sd-303, 8'sd-110}, {11'sd-982, 12'sd-1366, 11'sd-825}, {13'sd-2144, 12'sd1953, 13'sd2525}},
{{11'sd856, 13'sd2951, 13'sd3039}, {11'sd-809, 13'sd-2721, 13'sd2172}, {14'sd5299, 13'sd3244, 13'sd3719}},
{{8'sd-108, 12'sd1793, 13'sd-3625}, {12'sd1663, 13'sd-2906, 12'sd-1426}, {10'sd296, 10'sd-477, 7'sd37}},
{{11'sd640, 13'sd-2598, 12'sd1732}, {13'sd-2056, 13'sd2435, 13'sd2629}, {12'sd-1918, 10'sd-336, 12'sd1776}},
{{12'sd-1990, 13'sd2212, 11'sd-763}, {12'sd-2025, 12'sd1368, 12'sd1120}, {12'sd-1094, 12'sd1393, 12'sd1200}},
{{11'sd939, 12'sd1417, 10'sd-435}, {8'sd-112, 11'sd-986, 12'sd1545}, {12'sd-1777, 13'sd-2192, 9'sd-135}},
{{12'sd1698, 12'sd-1446, 8'sd-73}, {12'sd1853, 11'sd571, 13'sd-2252}, {8'sd69, 11'sd-1006, 12'sd-1599}},
{{11'sd700, 9'sd-158, 12'sd-1603}, {10'sd-473, 13'sd2968, 13'sd2170}, {13'sd3275, 12'sd1744, 11'sd-678}},
{{13'sd3431, 12'sd1735, 11'sd-760}, {13'sd2648, 13'sd2075, 13'sd-2943}, {12'sd1976, 12'sd-1206, 12'sd1651}},
{{11'sd914, 8'sd-87, 12'sd1953}, {12'sd-1443, 8'sd-81, 13'sd-2176}, {12'sd1701, 13'sd-4047, 12'sd-1767}},
{{13'sd-3819, 13'sd-2417, 11'sd547}, {13'sd-2987, 7'sd34, 13'sd2469}, {13'sd-3403, 14'sd-4182, 11'sd616}},
{{13'sd-2452, 13'sd-2302, 13'sd-2765}, {13'sd-2293, 9'sd140, 13'sd2640}, {11'sd-875, 13'sd-3031, 14'sd-4151}},
{{11'sd-1013, 12'sd1899, 12'sd1745}, {10'sd-378, 12'sd1358, 12'sd1168}, {10'sd-266, 12'sd-1065, 13'sd-2508}},
{{10'sd-478, 12'sd1580, 11'sd-652}, {11'sd-749, 12'sd1439, 12'sd1423}, {9'sd-249, 12'sd1117, 11'sd-840}},
{{13'sd-2456, 11'sd548, 12'sd-1132}, {12'sd-1877, 12'sd1057, 12'sd-1975}, {13'sd-2770, 12'sd-1489, 13'sd2223}},
{{12'sd1352, 13'sd2393, 13'sd-2692}, {11'sd986, 11'sd988, 12'sd-1194}, {13'sd-3141, 7'sd54, 10'sd270}},
{{12'sd-1428, 13'sd-3662, 13'sd-3145}, {11'sd-783, 12'sd-1500, 8'sd125}, {11'sd-619, 12'sd1277, 11'sd570}},
{{13'sd-3267, 8'sd-71, 10'sd420}, {12'sd1396, 11'sd-906, 8'sd-79}, {13'sd-2325, 12'sd1938, 11'sd679}},
{{13'sd3367, 10'sd474, 14'sd4424}, {14'sd4103, 11'sd-905, 13'sd2662}, {13'sd2864, 13'sd3182, 13'sd2985}},
{{12'sd-1758, 11'sd823, 12'sd-1396}, {11'sd622, 12'sd-1175, 12'sd-1477}, {13'sd2481, 10'sd281, 11'sd-588}},
{{11'sd-568, 9'sd-163, 11'sd1008}, {12'sd-1760, 7'sd34, 12'sd1809}, {13'sd2229, 12'sd1695, 12'sd-1529}},
{{13'sd2765, 10'sd-402, 10'sd275}, {4'sd4, 11'sd-673, 10'sd-425}, {9'sd-157, 11'sd-527, 12'sd-1218}},
{{13'sd3037, 13'sd2944, 13'sd2187}, {11'sd-759, 11'sd-733, 12'sd-1911}, {11'sd-699, 9'sd-173, 13'sd3576}},
{{13'sd-3191, 10'sd-502, 13'sd-2376}, {13'sd-2605, 12'sd1315, 13'sd2272}, {13'sd3069, 11'sd787, 13'sd2914}},
{{12'sd2004, 12'sd-1548, 10'sd501}, {12'sd2010, 12'sd-1343, 11'sd-557}, {13'sd-2292, 13'sd-2554, 13'sd-2817}},
{{12'sd-1970, 9'sd-254, 12'sd1471}, {13'sd-2416, 13'sd-2784, 9'sd243}, {13'sd2767, 13'sd-2606, 13'sd-3589}},
{{13'sd-3283, 13'sd-2293, 13'sd-2739}, {11'sd737, 13'sd2687, 12'sd1705}, {12'sd1288, 12'sd1183, 12'sd-1685}},
{{13'sd3267, 13'sd2602, 11'sd718}, {9'sd135, 13'sd-2094, 12'sd-1514}, {11'sd738, 10'sd-426, 13'sd2982}},
{{12'sd1509, 10'sd-258, 11'sd773}, {11'sd997, 13'sd2720, 13'sd-2669}, {13'sd-4093, 11'sd-648, 12'sd-1527}},
{{12'sd1057, 12'sd1808, 13'sd-2755}, {11'sd-818, 13'sd-2518, 11'sd-929}, {13'sd-2198, 11'sd-836, 13'sd-2461}},
{{11'sd-590, 10'sd374, 10'sd-472}, {10'sd-380, 12'sd1723, 6'sd-27}, {12'sd1163, 9'sd-147, 11'sd846}},
{{12'sd1598, 12'sd1232, 11'sd-733}, {9'sd237, 13'sd2307, 10'sd-380}, {12'sd1428, 12'sd-2042, 13'sd2538}},
{{11'sd-793, 10'sd263, 12'sd1860}, {12'sd-1485, 13'sd2173, 12'sd1662}, {13'sd2460, 12'sd1058, 11'sd630}}},
{
{{11'sd-761, 12'sd-1133, 12'sd1807}, {12'sd-1415, 12'sd1033, 12'sd-1425}, {9'sd234, 8'sd110, 12'sd-1224}},
{{11'sd1009, 12'sd1644, 13'sd2048}, {10'sd501, 13'sd-2514, 13'sd-2630}, {12'sd1730, 5'sd-11, 12'sd-2029}},
{{14'sd-4595, 12'sd-1681, 13'sd-4066}, {12'sd1861, 11'sd-838, 12'sd1319}, {11'sd633, 13'sd-3402, 13'sd-3460}},
{{12'sd-1086, 13'sd2661, 12'sd-1677}, {12'sd-1999, 13'sd3695, 9'sd-154}, {13'sd3796, 11'sd-659, 13'sd3381}},
{{12'sd-1155, 11'sd-903, 13'sd2846}, {11'sd744, 12'sd-1968, 13'sd3206}, {10'sd-325, 12'sd-1487, 13'sd3074}},
{{9'sd251, 12'sd-1640, 12'sd-1185}, {12'sd-1981, 9'sd-181, 12'sd-1432}, {13'sd2064, 12'sd-1814, 11'sd-613}},
{{12'sd2026, 13'sd3146, 13'sd3163}, {12'sd-1838, 11'sd692, 11'sd986}, {14'sd-5627, 11'sd591, 12'sd-1197}},
{{13'sd-2291, 13'sd-2592, 13'sd3302}, {12'sd-1401, 11'sd-853, 12'sd-1619}, {13'sd-3732, 13'sd-2445, 12'sd-1180}},
{{13'sd2769, 12'sd-1742, 13'sd3581}, {13'sd2209, 11'sd820, 10'sd-430}, {13'sd2779, 11'sd-534, 10'sd306}},
{{12'sd1079, 13'sd2354, 11'sd-939}, {13'sd2438, 11'sd-708, 13'sd-2747}, {8'sd68, 13'sd-2405, 12'sd1769}},
{{11'sd862, 12'sd1354, 13'sd2533}, {13'sd-2091, 10'sd416, 10'sd-391}, {13'sd-2208, 12'sd1362, 11'sd-793}},
{{13'sd2595, 13'sd2262, 12'sd-1740}, {4'sd-5, 11'sd644, 12'sd-1741}, {9'sd172, 11'sd-748, 13'sd-3790}},
{{13'sd2589, 11'sd-781, 12'sd1338}, {14'sd4522, 12'sd-1305, 13'sd3742}, {13'sd2173, 13'sd3042, 11'sd-534}},
{{11'sd688, 13'sd-2290, 12'sd-1408}, {13'sd2832, 13'sd-2579, 12'sd1192}, {13'sd2304, 13'sd2408, 13'sd2665}},
{{13'sd2115, 13'sd-2325, 12'sd-1319}, {12'sd1402, 12'sd-1215, 12'sd-1252}, {13'sd2424, 14'sd4174, 14'sd4350}},
{{12'sd1302, 11'sd-606, 12'sd1416}, {12'sd1450, 12'sd1644, 13'sd3214}, {11'sd-978, 10'sd367, 13'sd2481}},
{{13'sd-3405, 12'sd-1642, 11'sd-525}, {12'sd-1880, 11'sd806, 12'sd-1739}, {12'sd-1413, 13'sd-2697, 11'sd-933}},
{{13'sd-2768, 13'sd2281, 11'sd-848}, {11'sd802, 13'sd2539, 9'sd-218}, {13'sd2159, 12'sd-1101, 10'sd-449}},
{{11'sd-734, 13'sd2383, 13'sd3875}, {10'sd-373, 12'sd1618, 10'sd301}, {13'sd-3386, 12'sd1392, 12'sd1892}},
{{13'sd2776, 12'sd-1707, 13'sd2305}, {12'sd-1718, 10'sd262, 13'sd-2413}, {12'sd-1232, 11'sd-844, 10'sd318}},
{{14'sd-5883, 13'sd-2559, 11'sd981}, {12'sd-1549, 12'sd1036, 12'sd1093}, {11'sd-1008, 12'sd-1427, 5'sd11}},
{{10'sd-489, 12'sd1873, 12'sd1373}, {11'sd-639, 8'sd99, 10'sd-289}, {11'sd645, 11'sd-902, 10'sd299}},
{{9'sd242, 13'sd2259, 8'sd126}, {13'sd2969, 13'sd2685, 13'sd3206}, {11'sd708, 13'sd-2163, 12'sd-1545}},
{{12'sd1116, 13'sd-2188, 13'sd3122}, {12'sd1458, 13'sd-2364, 10'sd265}, {10'sd-420, 12'sd1677, 12'sd-1164}},
{{13'sd-2230, 10'sd475, 11'sd-754}, {11'sd-612, 8'sd83, 12'sd-1565}, {12'sd-1972, 11'sd-903, 13'sd2060}},
{{12'sd1966, 12'sd1995, 10'sd-280}, {11'sd573, 12'sd-1711, 11'sd845}, {11'sd754, 10'sd492, 13'sd-2674}},
{{12'sd1396, 12'sd1624, 12'sd1488}, {12'sd-1851, 7'sd-47, 13'sd3287}, {12'sd-1593, 8'sd-68, 12'sd-1855}},
{{13'sd3940, 14'sd4746, 10'sd401}, {12'sd1812, 13'sd2464, 12'sd1848}, {13'sd-2251, 12'sd1422, 13'sd-2429}},
{{12'sd-1956, 11'sd-881, 13'sd3379}, {11'sd980, 8'sd-122, 12'sd1680}, {13'sd-2097, 13'sd2200, 10'sd466}},
{{13'sd3483, 12'sd-1362, 9'sd-205}, {13'sd-2177, 12'sd1056, 12'sd-1223}, {13'sd-2460, 12'sd-1523, 11'sd-828}},
{{6'sd16, 12'sd-1050, 7'sd62}, {13'sd-3211, 13'sd-2507, 12'sd1120}, {13'sd-2928, 13'sd-2322, 13'sd-3286}},
{{12'sd-1839, 12'sd1509, 12'sd1799}, {12'sd-1753, 8'sd-103, 13'sd2489}, {12'sd1830, 9'sd212, 13'sd2910}},
{{13'sd3508, 13'sd2748, 12'sd1791}, {12'sd-1717, 6'sd-24, 11'sd804}, {10'sd-295, 13'sd3338, 13'sd3882}},
{{12'sd-2040, 12'sd1224, 13'sd-2936}, {10'sd-299, 12'sd-1795, 3'sd2}, {12'sd-1035, 12'sd-1316, 12'sd-1295}},
{{13'sd2657, 12'sd2016, 11'sd765}, {11'sd822, 12'sd1770, 12'sd1853}, {13'sd-3859, 10'sd488, 12'sd1821}},
{{11'sd993, 10'sd-412, 9'sd136}, {13'sd2981, 13'sd3320, 12'sd1827}, {12'sd1055, 13'sd3156, 13'sd-2863}},
{{13'sd-2822, 11'sd-925, 13'sd3080}, {12'sd1053, 13'sd-3288, 12'sd-1247}, {12'sd1941, 13'sd2628, 12'sd1495}},
{{13'sd2256, 11'sd-589, 12'sd-2021}, {12'sd1127, 13'sd-2268, 12'sd-1740}, {12'sd-1370, 11'sd-963, 9'sd-139}},
{{12'sd1221, 11'sd-641, 10'sd-381}, {13'sd3276, 12'sd1843, 12'sd-1799}, {12'sd1830, 13'sd3182, 12'sd-1052}},
{{11'sd-541, 10'sd464, 13'sd2481}, {13'sd-2216, 11'sd803, 13'sd-2403}, {13'sd2927, 11'sd926, 13'sd2456}},
{{9'sd-215, 13'sd-2329, 14'sd4220}, {13'sd3492, 13'sd-3654, 12'sd-1158}, {12'sd1598, 11'sd-755, 9'sd146}},
{{10'sd281, 10'sd342, 9'sd-147}, {6'sd17, 11'sd-594, 12'sd-1771}, {3'sd-2, 13'sd-3677, 13'sd-2924}},
{{11'sd524, 11'sd608, 8'sd-91}, {11'sd548, 11'sd-697, 13'sd2260}, {9'sd171, 12'sd-1039, 12'sd1133}},
{{12'sd-1925, 11'sd932, 10'sd278}, {10'sd317, 10'sd404, 12'sd-2017}, {12'sd1780, 12'sd-1751, 12'sd2036}},
{{13'sd-3277, 10'sd423, 13'sd-2677}, {12'sd-1188, 11'sd-987, 12'sd-1822}, {11'sd646, 12'sd1698, 11'sd-710}},
{{12'sd-1252, 13'sd2230, 8'sd-67}, {12'sd-1715, 12'sd1216, 13'sd2190}, {12'sd-1792, 11'sd898, 10'sd-460}},
{{13'sd-2641, 12'sd-1953, 12'sd-1978}, {13'sd2788, 12'sd1319, 12'sd1302}, {12'sd-1653, 11'sd974, 13'sd-3104}},
{{12'sd-1597, 13'sd-2569, 13'sd2512}, {9'sd-233, 12'sd1966, 12'sd-1486}, {7'sd41, 12'sd-1836, 12'sd1042}},
{{14'sd-6857, 12'sd-1598, 13'sd2869}, {12'sd-1539, 10'sd-447, 11'sd-911}, {12'sd-1557, 12'sd1784, 13'sd3957}},
{{12'sd1216, 13'sd2214, 12'sd1587}, {13'sd2192, 13'sd2617, 13'sd3471}, {13'sd3862, 12'sd1659, 13'sd3258}},
{{13'sd-2173, 9'sd-147, 13'sd3882}, {12'sd-1878, 13'sd3225, 11'sd-664}, {11'sd799, 13'sd2351, 12'sd-1264}},
{{12'sd-1029, 12'sd1791, 10'sd-356}, {12'sd1587, 13'sd2429, 13'sd-2389}, {12'sd-1525, 8'sd72, 13'sd-2414}},
{{13'sd2820, 13'sd2964, 13'sd-3167}, {12'sd-1525, 12'sd-1132, 11'sd-791}, {12'sd-1911, 13'sd-2179, 12'sd-1998}},
{{9'sd195, 8'sd97, 13'sd3276}, {13'sd-3194, 11'sd-657, 13'sd2672}, {14'sd-4480, 10'sd325, 12'sd-1413}},
{{12'sd-1448, 12'sd-1142, 13'sd-4040}, {11'sd-577, 13'sd-2116, 13'sd-2544}, {12'sd1234, 12'sd1201, 13'sd-2183}},
{{12'sd-1618, 13'sd-2572, 12'sd1959}, {11'sd543, 13'sd-2273, 12'sd1569}, {12'sd1703, 11'sd-1023, 10'sd-445}},
{{13'sd3170, 12'sd-1308, 13'sd2276}, {13'sd3148, 12'sd-1595, 13'sd-3125}, {12'sd1652, 12'sd1534, 11'sd-627}},
{{13'sd2249, 13'sd2305, 13'sd2141}, {13'sd2778, 13'sd3319, 13'sd2461}, {11'sd-522, 12'sd-1301, 14'sd4840}},
{{11'sd-785, 12'sd1983, 12'sd1038}, {12'sd-1224, 10'sd-339, 10'sd-368}, {10'sd-375, 12'sd-1254, 11'sd-706}},
{{10'sd-284, 11'sd-610, 12'sd-1845}, {8'sd75, 9'sd210, 14'sd-4252}, {12'sd-1245, 11'sd538, 14'sd-4813}},
{{12'sd-1841, 12'sd1978, 11'sd757}, {12'sd1032, 12'sd-1589, 13'sd2481}, {11'sd612, 11'sd-525, 13'sd-2349}},
{{12'sd1379, 12'sd-1709, 14'sd4109}, {12'sd1372, 13'sd-2134, 9'sd-253}, {10'sd455, 12'sd-1603, 11'sd-804}},
{{11'sd588, 12'sd-1325, 11'sd-658}, {11'sd-544, 13'sd2583, 12'sd-1733}, {12'sd1748, 12'sd-1122, 12'sd-1724}},
{{13'sd-3693, 14'sd-4138, 10'sd-488}, {13'sd-2855, 12'sd1108, 12'sd1877}, {13'sd-2633, 13'sd-2062, 11'sd-554}}},
{
{{12'sd-1968, 11'sd-519, 13'sd2463}, {11'sd-858, 11'sd965, 11'sd928}, {11'sd-828, 9'sd-155, 11'sd904}},
{{13'sd-2569, 12'sd1696, 10'sd-271}, {12'sd-2043, 5'sd12, 12'sd1242}, {11'sd-524, 11'sd804, 12'sd-1864}},
{{12'sd-1727, 8'sd-93, 6'sd-29}, {11'sd-838, 13'sd-2515, 11'sd-606}, {11'sd560, 12'sd-1155, 13'sd-2650}},
{{13'sd-2604, 13'sd-3425, 12'sd1468}, {10'sd-471, 12'sd-1106, 11'sd-840}, {13'sd-2290, 12'sd-1568, 12'sd-2035}},
{{12'sd1702, 11'sd966, 9'sd235}, {13'sd2136, 12'sd2013, 11'sd-746}, {12'sd1987, 13'sd2950, 13'sd-2297}},
{{10'sd-500, 13'sd2048, 10'sd-371}, {13'sd-2506, 12'sd-1519, 13'sd-2466}, {12'sd1199, 13'sd-2158, 5'sd-8}},
{{12'sd-1323, 13'sd2524, 12'sd-1386}, {13'sd-3194, 13'sd2307, 8'sd103}, {14'sd4291, 14'sd4579, 12'sd1117}},
{{11'sd-916, 11'sd554, 11'sd-962}, {13'sd2312, 12'sd1473, 13'sd2233}, {14'sd5071, 14'sd4208, 8'sd-85}},
{{13'sd2296, 10'sd-491, 11'sd-896}, {14'sd-4096, 11'sd714, 9'sd-154}, {13'sd-2620, 12'sd1030, 13'sd3003}},
{{11'sd749, 10'sd-297, 13'sd-2432}, {12'sd1538, 12'sd1916, 11'sd-932}, {13'sd-2083, 13'sd2488, 12'sd-1421}},
{{12'sd1560, 12'sd-1986, 12'sd-1914}, {13'sd-3061, 13'sd-3154, 12'sd-2013}, {12'sd1687, 11'sd-1004, 12'sd1079}},
{{9'sd241, 13'sd2678, 13'sd2341}, {13'sd-3657, 9'sd233, 12'sd-1715}, {10'sd-320, 13'sd2393, 10'sd418}},
{{14'sd-5618, 7'sd37, 11'sd-811}, {13'sd-2983, 14'sd-5597, 10'sd-456}, {12'sd-1186, 12'sd-1744, 13'sd2736}},
{{12'sd-1836, 8'sd72, 10'sd-470}, {13'sd-3022, 12'sd-1418, 9'sd-133}, {13'sd2200, 13'sd2096, 12'sd1845}},
{{11'sd602, 10'sd-293, 12'sd1198}, {9'sd248, 12'sd1306, 13'sd3269}, {13'sd-3185, 12'sd1818, 12'sd1389}},
{{6'sd22, 9'sd-232, 13'sd2252}, {12'sd-1453, 12'sd1191, 13'sd2050}, {11'sd-711, 10'sd346, 12'sd-1401}},
{{11'sd681, 9'sd-224, 12'sd-1573}, {12'sd1920, 8'sd-121, 12'sd-2027}, {10'sd-315, 13'sd2386, 3'sd2}},
{{13'sd3829, 12'sd-1568, 12'sd-1798}, {13'sd2633, 13'sd-3993, 11'sd849}, {13'sd3503, 11'sd973, 11'sd574}},
{{11'sd-933, 11'sd681, 13'sd2632}, {9'sd-173, 13'sd3069, 10'sd472}, {9'sd182, 13'sd2820, 10'sd-296}},
{{13'sd2341, 11'sd-882, 9'sd-243}, {13'sd-2868, 9'sd204, 11'sd531}, {13'sd2291, 11'sd-772, 13'sd-2243}},
{{12'sd-1208, 12'sd-1280, 12'sd-1136}, {11'sd-967, 9'sd-172, 11'sd899}, {12'sd1628, 9'sd-171, 7'sd-56}},
{{12'sd-1190, 13'sd-2491, 12'sd-1452}, {12'sd-1545, 13'sd-2553, 13'sd2440}, {7'sd-45, 13'sd2181, 13'sd3059}},
{{10'sd-338, 11'sd767, 12'sd-1362}, {13'sd2952, 12'sd1582, 13'sd3196}, {11'sd-1021, 13'sd2264, 10'sd-391}},
{{12'sd-1129, 10'sd416, 10'sd315}, {13'sd2927, 12'sd-1220, 11'sd658}, {10'sd-483, 10'sd317, 12'sd1387}},
{{11'sd-787, 11'sd836, 12'sd-1279}, {13'sd-2329, 12'sd-1951, 11'sd-822}, {12'sd-1112, 12'sd-2043, 12'sd1918}},
{{13'sd-2701, 9'sd-193, 9'sd-166}, {11'sd-866, 12'sd1557, 10'sd355}, {13'sd2195, 11'sd-1017, 12'sd1662}},
{{12'sd-1401, 13'sd2758, 10'sd295}, {12'sd-1186, 12'sd-1046, 12'sd-1421}, {13'sd2627, 5'sd9, 11'sd-947}},
{{13'sd-3444, 11'sd-778, 13'sd2606}, {11'sd-956, 9'sd160, 13'sd2710}, {11'sd-627, 12'sd-1707, 13'sd2210}},
{{11'sd-879, 12'sd-1188, 12'sd-1369}, {13'sd-2316, 13'sd-3736, 11'sd893}, {12'sd-1760, 12'sd-1059, 12'sd1127}},
{{12'sd-1718, 13'sd2266, 12'sd1343}, {11'sd-816, 13'sd-2458, 13'sd-2112}, {12'sd1059, 13'sd-2456, 13'sd2841}},
{{13'sd-2688, 11'sd-923, 13'sd-2346}, {9'sd190, 4'sd-7, 12'sd-1523}, {10'sd366, 11'sd-946, 13'sd-3927}},
{{13'sd2555, 13'sd3088, 12'sd1731}, {12'sd-1161, 13'sd2699, 12'sd1106}, {11'sd-759, 11'sd-641, 12'sd-1030}},
{{12'sd1103, 11'sd-647, 10'sd292}, {11'sd-524, 12'sd-1668, 13'sd2164}, {10'sd-432, 12'sd1310, 10'sd440}},
{{12'sd-1706, 9'sd135, 12'sd-1931}, {13'sd-2447, 12'sd-1910, 14'sd-4514}, {5'sd13, 11'sd-816, 11'sd911}},
{{12'sd-2003, 11'sd807, 13'sd3977}, {10'sd383, 12'sd1281, 13'sd2543}, {8'sd76, 12'sd1119, 12'sd2007}},
{{12'sd1046, 13'sd-3170, 12'sd-1455}, {13'sd-3174, 12'sd-1830, 13'sd-2170}, {12'sd-1548, 11'sd-832, 4'sd-4}},
{{4'sd-5, 11'sd-887, 12'sd1270}, {12'sd-1798, 10'sd-336, 13'sd-3198}, {12'sd-1809, 12'sd-1292, 9'sd156}},
{{9'sd-233, 5'sd10, 13'sd2400}, {12'sd-1383, 12'sd-1091, 13'sd-3161}, {13'sd-2137, 12'sd-1611, 13'sd2292}},
{{12'sd-1098, 13'sd2458, 13'sd2266}, {13'sd-2867, 10'sd421, 13'sd2495}, {8'sd-79, 12'sd-1461, 12'sd1815}},
{{11'sd-609, 13'sd2423, 13'sd-2459}, {12'sd-1683, 13'sd2724, 12'sd-1030}, {13'sd-2788, 13'sd-2305, 12'sd-1805}},
{{13'sd2663, 11'sd879, 12'sd1167}, {13'sd2077, 14'sd4387, 12'sd1277}, {10'sd-395, 12'sd-1128, 11'sd669}},
{{12'sd1500, 13'sd2558, 9'sd-214}, {13'sd-2366, 11'sd768, 11'sd745}, {11'sd1001, 12'sd-1297, 11'sd597}},
{{11'sd-819, 12'sd1208, 11'sd598}, {13'sd-3962, 11'sd625, 13'sd2074}, {11'sd-588, 12'sd-1354, 11'sd875}},
{{11'sd518, 12'sd1795, 10'sd-281}, {9'sd-160, 12'sd1835, 13'sd-2710}, {12'sd-1177, 12'sd-1301, 12'sd-1270}},
{{12'sd-1219, 11'sd663, 8'sd-121}, {12'sd1039, 12'sd1387, 10'sd-488}, {12'sd-1346, 13'sd3654, 13'sd2501}},
{{12'sd1981, 12'sd1970, 12'sd1566}, {11'sd-913, 13'sd-3506, 12'sd1898}, {12'sd1741, 11'sd875, 13'sd-2667}},
{{12'sd-1162, 12'sd1846, 12'sd1958}, {12'sd1808, 13'sd-3271, 12'sd-1931}, {13'sd-2166, 12'sd1552, 12'sd1787}},
{{13'sd3303, 13'sd2714, 12'sd1678}, {11'sd-964, 13'sd-2250, 12'sd-1605}, {11'sd980, 13'sd-2228, 8'sd85}},
{{12'sd1046, 12'sd-2032, 9'sd165}, {12'sd1124, 13'sd3004, 13'sd-2615}, {14'sd4682, 8'sd80, 13'sd-3064}},
{{14'sd4987, 13'sd2640, 14'sd4380}, {11'sd739, 12'sd1448, 14'sd4806}, {10'sd-373, 12'sd-1314, 10'sd486}},
{{13'sd-2467, 14'sd4525, 13'sd4016}, {10'sd511, 14'sd4541, 14'sd5969}, {10'sd-311, 11'sd594, 13'sd2475}},
{{9'sd190, 11'sd-593, 13'sd-2307}, {11'sd-827, 13'sd2683, 9'sd132}, {13'sd-3709, 11'sd-739, 12'sd1864}},
{{12'sd-1631, 12'sd-1885, 11'sd-540}, {12'sd1714, 11'sd804, 13'sd2661}, {12'sd1680, 13'sd-2642, 13'sd2264}},
{{11'sd790, 11'sd870, 11'sd1007}, {11'sd945, 12'sd-1735, 12'sd1957}, {12'sd1561, 12'sd-1801, 12'sd-1838}},
{{9'sd-248, 10'sd385, 12'sd1642}, {12'sd-1786, 13'sd-3400, 12'sd1183}, {13'sd-2224, 12'sd-1530, 11'sd-568}},
{{11'sd-776, 11'sd-934, 10'sd-470}, {11'sd-815, 8'sd-92, 12'sd-1178}, {10'sd376, 9'sd-177, 9'sd187}},
{{14'sd-4348, 13'sd2985, 13'sd2202}, {13'sd-3584, 13'sd-2463, 11'sd-617}, {14'sd-5170, 11'sd-977, 12'sd1236}},
{{13'sd-4022, 13'sd-2934, 12'sd1595}, {10'sd-487, 13'sd-2163, 12'sd-1288}, {12'sd1419, 12'sd1884, 13'sd2300}},
{{13'sd-2615, 13'sd-3275, 14'sd-4453}, {12'sd-1681, 9'sd-143, 13'sd-3551}, {13'sd2521, 12'sd1941, 12'sd1131}},
{{10'sd-287, 13'sd-3408, 13'sd2660}, {13'sd-3694, 13'sd-3144, 11'sd-705}, {13'sd-3347, 12'sd-1945, 12'sd1062}},
{{12'sd-1499, 12'sd1565, 10'sd-407}, {13'sd3585, 13'sd3180, 11'sd-991}, {11'sd-883, 12'sd-1503, 12'sd1277}},
{{12'sd-1771, 12'sd-1100, 12'sd1396}, {13'sd2888, 13'sd2736, 8'sd-116}, {13'sd3946, 12'sd-1749, 12'sd-1685}},
{{14'sd-4291, 12'sd-1149, 12'sd1466}, {10'sd-268, 12'sd1872, 13'sd3337}, {13'sd-2064, 12'sd1637, 12'sd1713}},
{{13'sd2119, 11'sd-518, 9'sd-232}, {13'sd3497, 12'sd1761, 8'sd112}, {12'sd1754, 13'sd3236, 9'sd-128}}},
{
{{12'sd-1045, 12'sd-1214, 11'sd866}, {13'sd-2199, 13'sd-2631, 12'sd-1080}, {13'sd-3204, 13'sd-2645, 12'sd1411}},
{{12'sd1687, 10'sd-397, 13'sd2583}, {12'sd1284, 10'sd497, 12'sd-1069}, {11'sd-827, 12'sd-1698, 12'sd-1903}},
{{12'sd-1989, 12'sd-1458, 12'sd1719}, {11'sd882, 6'sd21, 12'sd1775}, {13'sd-3226, 14'sd-4715, 10'sd276}},
{{12'sd-1236, 12'sd1251, 12'sd1379}, {6'sd22, 10'sd280, 12'sd-1716}, {13'sd2616, 13'sd-2179, 11'sd828}},
{{13'sd-2631, 12'sd-1611, 13'sd2603}, {12'sd-1703, 11'sd-861, 12'sd-1937}, {11'sd-719, 4'sd5, 10'sd389}},
{{12'sd1512, 13'sd-2876, 12'sd-1687}, {11'sd906, 12'sd-1729, 12'sd-2029}, {13'sd2551, 13'sd2693, 12'sd-1046}},
{{12'sd1404, 9'sd237, 12'sd-1292}, {12'sd-2000, 13'sd-2982, 10'sd398}, {13'sd3539, 12'sd1665, 12'sd-1263}},
{{13'sd-3281, 11'sd-771, 12'sd-1248}, {11'sd708, 10'sd-382, 13'sd-2062}, {8'sd-127, 12'sd1615, 12'sd1168}},
{{13'sd2869, 12'sd1537, 13'sd-2166}, {11'sd-795, 13'sd-2522, 11'sd-908}, {12'sd1708, 12'sd1999, 11'sd-617}},
{{13'sd-2570, 12'sd1687, 9'sd177}, {12'sd1732, 5'sd-13, 8'sd-110}, {12'sd1888, 12'sd1235, 11'sd752}},
{{10'sd-440, 13'sd-2847, 12'sd-1721}, {11'sd-708, 9'sd-175, 12'sd-1979}, {9'sd-139, 12'sd1099, 13'sd-2434}},
{{12'sd-1186, 12'sd-1528, 12'sd-1271}, {12'sd1659, 11'sd-657, 12'sd-1706}, {11'sd-958, 6'sd26, 12'sd1477}},
{{13'sd-2726, 13'sd-3667, 12'sd-2002}, {13'sd-2764, 13'sd-3333, 12'sd-1957}, {11'sd889, 13'sd-3135, 13'sd2621}},
{{13'sd-2708, 12'sd-1361, 9'sd197}, {13'sd-2309, 11'sd527, 12'sd1399}, {10'sd-354, 12'sd-1428, 12'sd-1465}},
{{11'sd528, 12'sd-1242, 13'sd-2370}, {8'sd-71, 12'sd1545, 10'sd-511}, {13'sd-2172, 12'sd1793, 12'sd-1786}},
{{12'sd1910, 11'sd872, 13'sd2421}, {11'sd932, 12'sd1969, 13'sd-2220}, {11'sd992, 13'sd-2943, 7'sd-60}},
{{8'sd105, 13'sd-2281, 9'sd234}, {11'sd-833, 12'sd1133, 13'sd2734}, {13'sd2568, 9'sd242, 11'sd-706}},
{{11'sd-524, 12'sd1292, 13'sd2543}, {13'sd2824, 12'sd1912, 10'sd307}, {12'sd-1226, 12'sd1458, 12'sd2045}},
{{12'sd1529, 12'sd-1841, 11'sd1012}, {13'sd-2478, 12'sd1172, 11'sd1002}, {12'sd-1840, 11'sd-731, 12'sd-1513}},
{{11'sd-706, 11'sd-927, 12'sd1307}, {12'sd-1958, 13'sd-2844, 12'sd-1290}, {10'sd400, 11'sd588, 11'sd512}},
{{13'sd-3110, 10'sd497, 5'sd9}, {12'sd1435, 13'sd2207, 12'sd-1884}, {12'sd-1614, 12'sd1898, 13'sd-2251}},
{{11'sd857, 13'sd-3070, 12'sd1824}, {10'sd342, 13'sd-2955, 13'sd-2169}, {12'sd1551, 10'sd452, 12'sd-1639}},
{{12'sd-1922, 11'sd-945, 11'sd-726}, {12'sd1041, 12'sd1193, 12'sd1876}, {13'sd-2489, 12'sd1810, 12'sd1050}},
{{9'sd157, 12'sd-2013, 12'sd1846}, {13'sd2979, 11'sd777, 13'sd2775}, {12'sd-1236, 13'sd2659, 12'sd1129}},
{{10'sd341, 13'sd-2159, 11'sd-893}, {9'sd-230, 10'sd-482, 7'sd56}, {11'sd563, 12'sd1975, 11'sd668}},
{{12'sd-1050, 10'sd-441, 12'sd1323}, {11'sd979, 12'sd-1313, 11'sd669}, {12'sd1741, 11'sd662, 13'sd2161}},
{{12'sd-1915, 12'sd-1306, 11'sd1016}, {11'sd-602, 13'sd2680, 13'sd-2412}, {12'sd1705, 12'sd2031, 11'sd527}},
{{11'sd-691, 12'sd-1296, 12'sd1438}, {12'sd-1168, 11'sd673, 9'sd-226}, {11'sd-807, 13'sd2790, 11'sd844}},
{{12'sd-1749, 12'sd1567, 9'sd-232}, {13'sd-2689, 12'sd1362, 12'sd-1400}, {13'sd2219, 13'sd2681, 10'sd424}},
{{12'sd1435, 10'sd272, 11'sd-773}, {12'sd-1529, 12'sd1132, 11'sd585}, {13'sd2461, 11'sd-521, 11'sd806}},
{{11'sd-864, 13'sd3272, 11'sd926}, {12'sd-1054, 11'sd987, 12'sd1683}, {12'sd-1107, 13'sd2450, 12'sd-1906}},
{{12'sd1905, 11'sd-594, 12'sd-1471}, {12'sd1846, 13'sd2484, 10'sd487}, {12'sd1809, 13'sd2449, 11'sd-522}},
{{13'sd-2871, 9'sd-188, 12'sd1747}, {12'sd1261, 12'sd-1286, 13'sd2321}, {12'sd1251, 12'sd-1885, 10'sd-505}},
{{11'sd936, 11'sd-657, 13'sd-3972}, {12'sd1154, 13'sd-2486, 13'sd-2836}, {11'sd-649, 11'sd-541, 12'sd-1243}},
{{13'sd2719, 13'sd-2325, 8'sd74}, {13'sd2490, 12'sd-1374, 11'sd-615}, {13'sd-2373, 10'sd-389, 12'sd1883}},
{{13'sd2424, 13'sd-2728, 10'sd-491}, {13'sd-2623, 12'sd1932, 13'sd2423}, {10'sd-445, 12'sd1579, 10'sd495}},
{{10'sd-350, 9'sd-192, 10'sd-369}, {10'sd370, 12'sd-1491, 12'sd-1197}, {12'sd1880, 13'sd-2068, 11'sd601}},
{{11'sd937, 13'sd2747, 11'sd-867}, {10'sd328, 12'sd-2012, 13'sd-2386}, {9'sd173, 7'sd32, 9'sd-206}},
{{11'sd-970, 13'sd-2111, 4'sd-7}, {12'sd1630, 13'sd2401, 13'sd2287}, {12'sd-1720, 12'sd-1169, 13'sd-2479}},
{{12'sd1185, 13'sd2523, 13'sd-2726}, {13'sd-2631, 13'sd2594, 10'sd-456}, {13'sd-2166, 12'sd2047, 12'sd-1669}},
{{10'sd354, 13'sd-3028, 12'sd-1537}, {10'sd-461, 8'sd-101, 11'sd-514}, {12'sd1451, 13'sd-2536, 8'sd74}},
{{9'sd177, 11'sd-546, 12'sd-1771}, {13'sd-2109, 12'sd1788, 12'sd-1194}, {9'sd-207, 10'sd-335, 13'sd-2978}},
{{13'sd2765, 13'sd2371, 12'sd1555}, {10'sd301, 11'sd919, 11'sd-713}, {11'sd-907, 6'sd-21, 13'sd2831}},
{{13'sd-2083, 13'sd-2757, 12'sd-1579}, {12'sd-1953, 12'sd-1147, 12'sd1603}, {10'sd335, 13'sd-2807, 12'sd-1805}},
{{12'sd-1581, 12'sd-1712, 10'sd447}, {12'sd-1784, 8'sd81, 12'sd-1042}, {13'sd-2458, 12'sd1837, 11'sd840}},
{{13'sd2435, 12'sd-1176, 11'sd-628}, {12'sd1230, 12'sd1799, 11'sd691}, {12'sd1634, 12'sd-1320, 13'sd2103}},
{{12'sd1755, 13'sd-2511, 12'sd1927}, {12'sd1768, 12'sd-1528, 13'sd2609}, {12'sd-1770, 13'sd-2719, 12'sd-1289}},
{{10'sd-457, 13'sd-2835, 13'sd-3322}, {11'sd641, 11'sd-517, 13'sd-2589}, {7'sd-45, 12'sd-1216, 13'sd-2731}},
{{11'sd-832, 11'sd-552, 11'sd625}, {10'sd283, 12'sd-1236, 11'sd911}, {13'sd-2155, 13'sd3301, 13'sd3016}},
{{11'sd821, 12'sd-1685, 12'sd1471}, {12'sd-1874, 10'sd-344, 13'sd2651}, {9'sd-146, 13'sd-2607, 12'sd1707}},
{{10'sd377, 10'sd504, 13'sd3264}, {11'sd728, 12'sd-1034, 13'sd3320}, {12'sd-1943, 11'sd802, 13'sd2527}},
{{12'sd1273, 12'sd1670, 13'sd-2753}, {13'sd2411, 12'sd1470, 13'sd-3124}, {6'sd-22, 13'sd2161, 11'sd-702}},
{{12'sd-1570, 11'sd-953, 9'sd181}, {9'sd194, 13'sd-2301, 12'sd2022}, {11'sd682, 12'sd-1400, 10'sd-296}},
{{10'sd-364, 8'sd95, 12'sd-1360}, {6'sd18, 12'sd1071, 7'sd-38}, {12'sd1913, 12'sd-1252, 12'sd-1571}},
{{13'sd-2150, 10'sd481, 12'sd-1976}, {9'sd252, 8'sd83, 10'sd-411}, {9'sd-204, 13'sd-3043, 8'sd122}},
{{12'sd1168, 12'sd-1734, 10'sd-402}, {11'sd-860, 12'sd1491, 12'sd-1404}, {12'sd-1912, 13'sd2168, 11'sd-685}},
{{12'sd-1699, 12'sd-1386, 13'sd2332}, {13'sd-2347, 13'sd2523, 13'sd-2246}, {11'sd929, 13'sd-2134, 13'sd-2805}},
{{11'sd718, 13'sd2234, 12'sd1197}, {12'sd-1971, 9'sd179, 13'sd3205}, {12'sd1874, 12'sd1563, 11'sd981}},
{{8'sd-71, 12'sd1163, 10'sd-503}, {11'sd625, 11'sd-703, 7'sd-45}, {13'sd2136, 14'sd4115, 12'sd2018}},
{{11'sd553, 13'sd-2120, 11'sd-1019}, {12'sd-1674, 12'sd1261, 13'sd-2182}, {12'sd-1324, 11'sd746, 11'sd555}},
{{11'sd809, 10'sd304, 11'sd903}, {12'sd-1459, 13'sd-2071, 11'sd-774}, {12'sd-1275, 13'sd-2630, 7'sd-44}},
{{12'sd-1193, 12'sd-1291, 9'sd-248}, {11'sd635, 12'sd1264, 13'sd-2458}, {11'sd-1009, 7'sd56, 13'sd2427}},
{{11'sd-896, 11'sd-735, 12'sd1197}, {12'sd-1092, 12'sd-1639, 12'sd1051}, {13'sd-3893, 13'sd-2476, 13'sd2766}},
{{12'sd-2034, 10'sd323, 12'sd-1871}, {13'sd2106, 11'sd-586, 10'sd262}, {9'sd-223, 12'sd1548, 12'sd-1605}}},
{
{{13'sd2388, 13'sd2870, 12'sd-1024}, {12'sd1295, 13'sd-2344, 13'sd2590}, {8'sd107, 12'sd1754, 13'sd-2697}},
{{8'sd-74, 12'sd-1669, 12'sd-2016}, {9'sd-133, 10'sd-298, 11'sd-858}, {11'sd822, 11'sd-663, 11'sd911}},
{{14'sd5419, 10'sd314, 12'sd2035}, {11'sd-540, 10'sd397, 8'sd-100}, {10'sd-260, 12'sd-1680, 13'sd3081}},
{{12'sd1725, 13'sd2299, 12'sd1831}, {12'sd-1543, 10'sd438, 5'sd-13}, {13'sd2363, 13'sd-2184, 13'sd-2473}},
{{11'sd755, 10'sd-502, 12'sd-1280}, {12'sd-2029, 13'sd2753, 9'sd225}, {12'sd1954, 12'sd-2033, 12'sd1200}},
{{12'sd-1899, 12'sd-1272, 10'sd352}, {10'sd-379, 12'sd1686, 13'sd2586}, {11'sd-971, 12'sd-1285, 10'sd449}},
{{12'sd1237, 10'sd-291, 13'sd-3158}, {13'sd2282, 12'sd1296, 12'sd1630}, {14'sd4343, 13'sd2740, 12'sd-1297}},
{{13'sd3657, 13'sd2296, 13'sd2874}, {12'sd1945, 9'sd144, 13'sd3086}, {13'sd2659, 10'sd-442, 13'sd3462}},
{{13'sd-2184, 11'sd-703, 12'sd-1447}, {12'sd1041, 13'sd2110, 12'sd1790}, {13'sd-2784, 12'sd-1267, 12'sd-1076}},
{{11'sd574, 12'sd1689, 12'sd-1932}, {12'sd-1116, 12'sd-1045, 12'sd1790}, {11'sd866, 13'sd-2328, 13'sd2228}},
{{9'sd-197, 12'sd-1061, 12'sd2034}, {13'sd2149, 12'sd1194, 8'sd117}, {13'sd-2185, 13'sd-2597, 12'sd-1402}},
{{12'sd-1830, 12'sd-1285, 12'sd1301}, {12'sd-1964, 12'sd1454, 12'sd1102}, {12'sd-1093, 13'sd-2684, 12'sd1766}},
{{13'sd-2620, 12'sd1258, 12'sd-1437}, {13'sd-3818, 13'sd-2396, 12'sd1370}, {12'sd-1045, 13'sd3021, 9'sd245}},
{{13'sd-2124, 12'sd1675, 12'sd-1130}, {12'sd1781, 11'sd-762, 12'sd-1637}, {11'sd-515, 9'sd-190, 13'sd-2287}},
{{13'sd2438, 12'sd1208, 12'sd2044}, {7'sd-48, 11'sd-782, 13'sd-2901}, {11'sd-948, 8'sd74, 12'sd1549}},
{{8'sd-110, 13'sd-2212, 12'sd-1659}, {12'sd-1118, 12'sd-1698, 13'sd-2532}, {13'sd-2859, 12'sd-1818, 12'sd-1489}},
{{12'sd1284, 11'sd866, 12'sd-1530}, {8'sd-96, 12'sd-1475, 10'sd315}, {13'sd-2425, 9'sd175, 10'sd-329}},
{{14'sd-5691, 12'sd-1839, 11'sd-662}, {12'sd1368, 13'sd-2598, 9'sd179}, {12'sd1943, 12'sd1495, 9'sd-180}},
{{11'sd597, 11'sd-913, 10'sd420}, {12'sd-1395, 10'sd482, 12'sd1582}, {9'sd-149, 9'sd-224, 11'sd-857}},
{{12'sd-1326, 11'sd-551, 11'sd-622}, {11'sd-1023, 11'sd-801, 12'sd-1048}, {12'sd1220, 9'sd200, 12'sd1105}},
{{9'sd176, 12'sd1224, 12'sd1956}, {12'sd-1292, 12'sd1941, 11'sd741}, {12'sd-1651, 13'sd-2059, 14'sd-4477}},
{{12'sd1340, 8'sd121, 13'sd3051}, {13'sd-3016, 13'sd-2574, 13'sd-2326}, {7'sd45, 11'sd-994, 11'sd-776}},
{{13'sd3078, 13'sd-2060, 12'sd1503}, {12'sd-1998, 10'sd-475, 11'sd-888}, {12'sd-1801, 12'sd-1366, 11'sd-874}},
{{12'sd-1435, 13'sd-2343, 12'sd-1377}, {13'sd2396, 13'sd-2525, 12'sd1514}, {12'sd-1271, 12'sd1527, 13'sd-3020}},
{{13'sd2714, 10'sd-333, 9'sd146}, {11'sd553, 12'sd-1439, 11'sd-746}, {11'sd644, 12'sd1549, 13'sd2249}},
{{12'sd1039, 12'sd1191, 13'sd-2214}, {12'sd-1221, 11'sd852, 11'sd973}, {9'sd136, 12'sd1868, 12'sd-1958}},
{{12'sd-1818, 12'sd-1855, 11'sd-985}, {12'sd-1646, 9'sd232, 12'sd-1309}, {13'sd2872, 9'sd233, 13'sd2583}},
{{11'sd584, 12'sd1619, 13'sd-2095}, {8'sd-99, 13'sd3083, 10'sd286}, {13'sd3003, 13'sd2227, 13'sd3407}},
{{12'sd1400, 7'sd36, 10'sd265}, {12'sd1459, 12'sd-1796, 11'sd-870}, {9'sd134, 9'sd-233, 13'sd-2464}},
{{12'sd-1993, 12'sd-1140, 11'sd959}, {13'sd2253, 9'sd183, 13'sd2064}, {12'sd1343, 13'sd-2496, 8'sd-79}},
{{12'sd-1434, 14'sd-5643, 13'sd-2292}, {12'sd-1596, 12'sd-1442, 11'sd-599}, {14'sd4274, 11'sd740, 12'sd-1615}},
{{11'sd544, 12'sd-1506, 13'sd-2467}, {13'sd-2694, 11'sd728, 13'sd-2073}, {12'sd-1560, 11'sd-652, 13'sd2308}},
{{12'sd-1585, 12'sd-1883, 13'sd-2484}, {10'sd-391, 13'sd-3442, 11'sd-861}, {12'sd1419, 11'sd-893, 13'sd-3985}},
{{11'sd-558, 12'sd-1057, 14'sd4331}, {8'sd82, 11'sd-780, 12'sd1885}, {7'sd60, 13'sd2617, 13'sd3893}},
{{12'sd-1730, 12'sd1324, 13'sd-2788}, {13'sd3285, 11'sd-775, 13'sd2643}, {11'sd-729, 12'sd1320, 12'sd-1299}},
{{13'sd-2119, 13'sd2203, 12'sd2041}, {10'sd460, 13'sd-2682, 13'sd2169}, {12'sd1670, 10'sd-318, 11'sd1015}},
{{13'sd2514, 12'sd1294, 12'sd-1054}, {10'sd259, 11'sd900, 12'sd-1983}, {13'sd-2071, 12'sd1743, 12'sd1139}},
{{13'sd-2757, 11'sd-696, 13'sd-3036}, {11'sd-1012, 11'sd-810, 12'sd1622}, {13'sd2178, 13'sd-2072, 12'sd1781}},
{{12'sd-1580, 10'sd400, 13'sd2276}, {12'sd-1043, 10'sd506, 10'sd-266}, {12'sd1071, 12'sd-1279, 11'sd998}},
{{13'sd2053, 12'sd1869, 11'sd-612}, {11'sd862, 11'sd957, 11'sd907}, {12'sd1247, 11'sd-652, 12'sd-1842}},
{{12'sd-1648, 13'sd3668, 12'sd-1069}, {12'sd-1346, 13'sd2292, 13'sd-2163}, {13'sd-3271, 12'sd-1743, 8'sd108}},
{{13'sd2128, 11'sd642, 11'sd-720}, {11'sd963, 12'sd-1389, 12'sd-1275}, {9'sd148, 12'sd-1775, 11'sd-807}},
{{11'sd805, 11'sd-818, 13'sd-2561}, {13'sd-2598, 12'sd-1728, 11'sd-802}, {12'sd-1336, 12'sd-1242, 5'sd-11}},
{{12'sd-1358, 13'sd-2644, 12'sd-1950}, {12'sd-1653, 12'sd-1144, 13'sd-2952}, {12'sd1885, 13'sd2542, 13'sd2665}},
{{12'sd1796, 13'sd2097, 11'sd641}, {10'sd308, 10'sd412, 12'sd-1663}, {10'sd499, 10'sd293, 12'sd-2034}},
{{12'sd-1107, 13'sd2697, 12'sd1697}, {13'sd-2708, 11'sd668, 11'sd-878}, {13'sd-2101, 12'sd-1768, 11'sd-952}},
{{11'sd962, 12'sd1617, 13'sd2579}, {13'sd-2659, 13'sd-2372, 12'sd1047}, {11'sd866, 11'sd-920, 12'sd-1328}},
{{14'sd4276, 10'sd369, 12'sd-1520}, {10'sd-259, 13'sd-2470, 12'sd-1517}, {13'sd2200, 11'sd-901, 12'sd1321}},
{{13'sd-2088, 12'sd-1703, 13'sd-2936}, {13'sd3448, 12'sd1823, 11'sd-965}, {12'sd1452, 13'sd-2931, 11'sd807}},
{{13'sd-3901, 10'sd442, 13'sd-3582}, {13'sd-3139, 12'sd-1277, 11'sd-655}, {13'sd2566, 13'sd2243, 10'sd294}},
{{12'sd1159, 10'sd422, 8'sd-74}, {12'sd-1244, 11'sd-990, 11'sd-969}, {13'sd-2586, 11'sd-710, 13'sd2202}},
{{11'sd639, 12'sd1962, 13'sd-2415}, {10'sd505, 12'sd1875, 11'sd-574}, {12'sd1511, 12'sd1391, 9'sd150}},
{{13'sd-2134, 7'sd45, 13'sd2164}, {13'sd-2497, 10'sd281, 11'sd-806}, {13'sd2814, 10'sd463, 13'sd2574}},
{{11'sd-554, 13'sd2233, 10'sd-295}, {11'sd-936, 10'sd-461, 9'sd232}, {11'sd-841, 12'sd-1221, 12'sd-1521}},
{{12'sd-1267, 10'sd363, 8'sd-72}, {11'sd861, 13'sd-2109, 12'sd1499}, {12'sd1086, 12'sd-1360, 13'sd2872}},
{{12'sd1338, 12'sd1715, 13'sd-2308}, {12'sd-1199, 12'sd-1401, 12'sd-1317}, {9'sd-254, 12'sd-1141, 12'sd-1221}},
{{12'sd1956, 13'sd2536, 13'sd2458}, {11'sd-802, 4'sd-6, 12'sd-2043}, {13'sd-2915, 12'sd-1897, 13'sd2633}},
{{13'sd-2072, 11'sd795, 11'sd-722}, {10'sd-437, 13'sd2512, 8'sd117}, {12'sd1821, 12'sd1504, 12'sd1657}},
{{11'sd746, 10'sd-397, 11'sd-690}, {13'sd2576, 6'sd17, 13'sd-2546}, {12'sd1526, 11'sd-825, 12'sd-1595}},
{{9'sd-226, 9'sd202, 12'sd1466}, {12'sd-1331, 12'sd1336, 8'sd124}, {13'sd2624, 10'sd-259, 11'sd679}},
{{13'sd-2789, 13'sd-2833, 12'sd1220}, {13'sd2455, 12'sd-1993, 12'sd1364}, {12'sd-1138, 11'sd-679, 13'sd2837}},
{{12'sd1439, 11'sd819, 13'sd-2475}, {10'sd491, 12'sd-1717, 10'sd-473}, {10'sd-266, 9'sd-203, 13'sd2283}},
{{12'sd-1310, 10'sd382, 10'sd280}, {12'sd1274, 13'sd-2865, 13'sd-2172}, {11'sd833, 12'sd1218, 12'sd1665}},
{{11'sd819, 10'sd412, 13'sd-2092}, {12'sd-1456, 12'sd1740, 12'sd1990}, {13'sd2245, 13'sd2246, 13'sd-2079}}},
{
{{13'sd-2858, 11'sd-698, 9'sd-205}, {13'sd-2979, 13'sd2067, 9'sd183}, {12'sd1350, 12'sd1795, 12'sd2034}},
{{12'sd-1913, 13'sd-2925, 13'sd-2318}, {12'sd-1945, 10'sd360, 10'sd-422}, {12'sd1438, 12'sd-1105, 12'sd1639}},
{{13'sd-2204, 12'sd-1715, 13'sd-3957}, {12'sd-1468, 12'sd1683, 12'sd-2039}, {7'sd62, 10'sd299, 10'sd417}},
{{12'sd-1201, 10'sd-418, 12'sd-1391}, {12'sd1528, 13'sd2054, 13'sd-2378}, {11'sd-940, 10'sd507, 10'sd411}},
{{13'sd2070, 13'sd2258, 12'sd1337}, {12'sd1861, 10'sd360, 4'sd-5}, {11'sd872, 9'sd-157, 13'sd2739}},
{{13'sd-2882, 10'sd-500, 13'sd2914}, {11'sd714, 12'sd1867, 11'sd559}, {12'sd1775, 13'sd2315, 6'sd-26}},
{{6'sd-23, 11'sd630, 13'sd-3410}, {11'sd975, 12'sd1907, 12'sd1873}, {12'sd-1474, 11'sd773, 13'sd-3852}},
{{12'sd1989, 12'sd-1833, 10'sd-327}, {11'sd517, 11'sd-1023, 13'sd-2672}, {12'sd1878, 13'sd-3019, 11'sd-523}},
{{13'sd2408, 12'sd-1178, 13'sd2124}, {13'sd3282, 12'sd-2018, 12'sd-1039}, {12'sd-1190, 13'sd-2745, 12'sd1237}},
{{11'sd-890, 12'sd1519, 11'sd692}, {12'sd-1533, 12'sd1956, 12'sd-1413}, {11'sd789, 12'sd2028, 11'sd818}},
{{11'sd-873, 9'sd-183, 11'sd995}, {12'sd-1917, 12'sd-1241, 10'sd-321}, {12'sd1852, 12'sd-1304, 13'sd-2206}},
{{13'sd-2885, 11'sd-820, 12'sd-1430}, {13'sd-2178, 7'sd33, 11'sd872}, {10'sd-478, 11'sd-1009, 12'sd-1508}},
{{13'sd-3037, 13'sd2308, 13'sd-2415}, {12'sd-1061, 11'sd707, 8'sd-102}, {11'sd583, 13'sd2209, 12'sd-1380}},
{{12'sd-1544, 13'sd-2827, 12'sd1285}, {12'sd-1282, 13'sd2170, 12'sd-1294}, {12'sd-1387, 13'sd-2803, 10'sd-421}},
{{11'sd-616, 8'sd68, 11'sd-710}, {12'sd1741, 13'sd3046, 12'sd-1298}, {12'sd1952, 12'sd1060, 10'sd-358}},
{{12'sd1403, 13'sd2131, 13'sd-2812}, {13'sd-2573, 7'sd36, 10'sd403}, {12'sd-1608, 9'sd137, 12'sd-1949}},
{{12'sd-1807, 10'sd399, 11'sd-595}, {13'sd2393, 12'sd1532, 10'sd351}, {11'sd986, 8'sd-87, 10'sd-370}},
{{12'sd1760, 12'sd1196, 11'sd-761}, {13'sd3118, 11'sd-803, 11'sd-712}, {13'sd3031, 13'sd2612, 11'sd781}},
{{13'sd2638, 12'sd1324, 12'sd-1794}, {12'sd-1620, 13'sd-2058, 8'sd116}, {12'sd1389, 13'sd2083, 11'sd-1002}},
{{12'sd1724, 12'sd1222, 12'sd1098}, {9'sd142, 11'sd1010, 11'sd614}, {11'sd-746, 13'sd2137, 12'sd1778}},
{{8'sd-87, 13'sd2067, 11'sd-852}, {11'sd-580, 13'sd2229, 10'sd486}, {12'sd-1916, 12'sd-1156, 12'sd1562}},
{{13'sd2964, 9'sd208, 12'sd1346}, {13'sd3119, 13'sd2782, 11'sd-580}, {10'sd-459, 13'sd2957, 11'sd-920}},
{{9'sd-193, 12'sd-1451, 13'sd2702}, {12'sd1775, 12'sd-1559, 13'sd2061}, {11'sd903, 12'sd1219, 11'sd731}},
{{12'sd1814, 12'sd-1664, 11'sd-618}, {12'sd-1029, 11'sd-894, 12'sd-1972}, {12'sd-1281, 11'sd920, 11'sd-955}},
{{13'sd-2186, 11'sd867, 12'sd1895}, {12'sd1911, 10'sd377, 12'sd2044}, {13'sd-2092, 12'sd-1691, 9'sd172}},
{{13'sd-2118, 12'sd1388, 13'sd-2387}, {13'sd-2427, 10'sd283, 12'sd1948}, {12'sd1251, 11'sd567, 13'sd2108}},
{{13'sd-2805, 12'sd-1383, 12'sd-1280}, {12'sd-1749, 11'sd784, 13'sd-2266}, {11'sd-534, 9'sd183, 11'sd-752}},
{{13'sd2867, 12'sd1585, 13'sd3702}, {12'sd-1787, 11'sd-819, 11'sd789}, {12'sd-2000, 11'sd-1009, 10'sd-475}},
{{12'sd1616, 12'sd1378, 11'sd-965}, {12'sd1073, 12'sd-1205, 12'sd-1158}, {12'sd-1962, 12'sd-2007, 10'sd471}},
{{11'sd-914, 12'sd1243, 13'sd-2715}, {13'sd-2211, 8'sd-118, 13'sd2671}, {11'sd-673, 12'sd1540, 13'sd2424}},
{{13'sd3613, 8'sd-64, 10'sd312}, {13'sd3667, 13'sd3544, 13'sd3508}, {13'sd2794, 10'sd-283, 14'sd4414}},
{{12'sd1921, 11'sd765, 12'sd1314}, {13'sd2445, 12'sd-1259, 12'sd1857}, {12'sd1706, 13'sd2391, 7'sd-33}},
{{13'sd-2223, 7'sd32, 13'sd3121}, {12'sd-1897, 12'sd1914, 12'sd1572}, {13'sd-3477, 12'sd-1404, 12'sd-1399}},
{{13'sd-2776, 12'sd1568, 13'sd-2215}, {10'sd271, 13'sd-2467, 11'sd866}, {12'sd1551, 12'sd-1742, 12'sd1309}},
{{12'sd1796, 10'sd462, 13'sd2432}, {12'sd-1071, 12'sd-1338, 13'sd2384}, {12'sd-1634, 12'sd1462, 13'sd2048}},
{{13'sd2446, 9'sd193, 13'sd-2163}, {12'sd-1985, 12'sd-1105, 10'sd-357}, {13'sd-2239, 13'sd-2215, 11'sd632}},
{{12'sd1467, 12'sd1872, 13'sd2754}, {13'sd2205, 13'sd-2800, 13'sd-2484}, {12'sd1239, 13'sd-2200, 12'sd1821}},
{{12'sd1726, 11'sd996, 13'sd-2186}, {9'sd132, 13'sd-2517, 11'sd679}, {12'sd1172, 11'sd554, 12'sd1415}},
{{13'sd-3866, 12'sd-1726, 12'sd1209}, {11'sd-717, 10'sd-260, 11'sd-840}, {13'sd-3969, 13'sd-2387, 12'sd1261}},
{{7'sd-50, 11'sd828, 11'sd848}, {11'sd658, 9'sd227, 10'sd385}, {12'sd-1246, 13'sd-2290, 11'sd-929}},
{{11'sd698, 9'sd-158, 13'sd-2093}, {13'sd3273, 12'sd-1510, 12'sd-1399}, {10'sd386, 12'sd-1288, 10'sd-474}},
{{14'sd-4270, 13'sd-3521, 12'sd1365}, {13'sd-2791, 13'sd-2710, 12'sd1402}, {13'sd3488, 13'sd3808, 13'sd2807}},
{{11'sd-909, 12'sd-1731, 12'sd-1953}, {11'sd848, 12'sd1709, 12'sd-1540}, {12'sd-1420, 12'sd1671, 12'sd1914}},
{{12'sd1274, 11'sd689, 13'sd2464}, {12'sd1613, 12'sd-1868, 13'sd2319}, {12'sd-1471, 13'sd2302, 12'sd1338}},
{{12'sd-1737, 11'sd-661, 9'sd181}, {11'sd767, 13'sd2079, 11'sd691}, {12'sd-1335, 10'sd508, 12'sd-1935}},
{{12'sd1723, 10'sd495, 11'sd-848}, {13'sd2753, 12'sd-1392, 11'sd692}, {11'sd-702, 13'sd-2291, 12'sd1799}},
{{13'sd2100, 9'sd-223, 13'sd2177}, {12'sd1394, 11'sd635, 9'sd-242}, {12'sd-1039, 11'sd-961, 11'sd731}},
{{9'sd-131, 13'sd-2451, 13'sd-2714}, {11'sd581, 11'sd-983, 10'sd393}, {11'sd-937, 11'sd-937, 12'sd1184}},
{{12'sd1688, 10'sd455, 13'sd-2869}, {11'sd-523, 12'sd-1671, 13'sd-2517}, {13'sd2168, 10'sd467, 12'sd-1606}},
{{13'sd3420, 11'sd-878, 12'sd1635}, {11'sd940, 10'sd502, 12'sd1136}, {9'sd189, 12'sd1271, 11'sd-1014}},
{{10'sd-420, 13'sd-2224, 10'sd259}, {12'sd-1130, 13'sd-2976, 12'sd1129}, {10'sd-296, 13'sd3396, 11'sd786}},
{{7'sd53, 9'sd-250, 12'sd2021}, {11'sd999, 9'sd-249, 8'sd-66}, {11'sd1013, 10'sd306, 12'sd1440}},
{{12'sd-1892, 13'sd2586, 11'sd-813}, {12'sd-1853, 10'sd-293, 11'sd-547}, {10'sd414, 12'sd-1447, 10'sd396}},
{{10'sd-338, 12'sd1545, 10'sd-373}, {13'sd2725, 13'sd-2749, 13'sd-2253}, {11'sd-549, 9'sd175, 12'sd-1244}},
{{13'sd-2903, 12'sd2016, 12'sd-1904}, {13'sd-3518, 11'sd595, 12'sd-1351}, {13'sd-2129, 10'sd433, 12'sd1224}},
{{13'sd2488, 12'sd1527, 13'sd-2340}, {11'sd901, 12'sd1785, 10'sd-439}, {11'sd-562, 13'sd2169, 11'sd-829}},
{{10'sd-406, 11'sd943, 12'sd-1983}, {13'sd-3158, 12'sd-1142, 11'sd796}, {11'sd755, 12'sd-1990, 13'sd2682}},
{{11'sd-885, 13'sd2669, 13'sd-2445}, {10'sd404, 12'sd1390, 12'sd-1698}, {11'sd786, 12'sd-1709, 13'sd-2791}},
{{13'sd-3586, 11'sd891, 9'sd255}, {13'sd-3539, 10'sd338, 9'sd-232}, {11'sd-805, 10'sd-299, 13'sd-3553}},
{{12'sd-1978, 11'sd773, 12'sd1232}, {10'sd-313, 12'sd1594, 11'sd619}, {10'sd-378, 12'sd-1125, 12'sd-1559}},
{{12'sd1315, 13'sd2687, 11'sd877}, {11'sd-671, 9'sd-128, 12'sd1373}, {5'sd15, 9'sd-208, 12'sd1382}},
{{13'sd2054, 11'sd775, 12'sd1846}, {12'sd-1164, 13'sd2103, 12'sd1354}, {13'sd-2897, 12'sd1261, 12'sd-1526}},
{{13'sd-2726, 11'sd631, 10'sd420}, {13'sd-2048, 11'sd896, 12'sd-1242}, {10'sd-297, 11'sd936, 12'sd-1339}},
{{13'sd-2451, 10'sd-317, 13'sd-2197}, {13'sd2385, 12'sd-1293, 12'sd-1757}, {12'sd1526, 11'sd656, 13'sd2606}}},
{
{{13'sd-2832, 12'sd-2012, 12'sd1658}, {10'sd-438, 12'sd-1385, 10'sd489}, {13'sd-2785, 11'sd714, 12'sd-1783}},
{{9'sd-166, 13'sd-2297, 11'sd-655}, {11'sd652, 12'sd1351, 13'sd-2504}, {11'sd844, 13'sd2620, 11'sd993}},
{{12'sd-2035, 10'sd328, 11'sd866}, {9'sd-154, 13'sd2698, 12'sd2033}, {13'sd-2947, 7'sd34, 12'sd-1170}},
{{11'sd870, 9'sd149, 11'sd661}, {11'sd-623, 12'sd1034, 12'sd-1775}, {13'sd-2373, 11'sd602, 12'sd1162}},
{{13'sd2907, 12'sd-2032, 11'sd-844}, {10'sd374, 13'sd2271, 13'sd-2467}, {13'sd2783, 13'sd2337, 12'sd1117}},
{{8'sd94, 12'sd1318, 13'sd2225}, {12'sd1025, 11'sd-602, 13'sd-2276}, {12'sd2018, 12'sd-1024, 10'sd-425}},
{{12'sd-1072, 12'sd2007, 11'sd955}, {11'sd952, 13'sd2721, 12'sd1130}, {11'sd-621, 13'sd3407, 6'sd24}},
{{13'sd-2133, 13'sd-3206, 13'sd-3626}, {9'sd-246, 13'sd-2502, 12'sd1154}, {11'sd888, 12'sd-1636, 13'sd-2503}},
{{12'sd-1076, 9'sd-177, 13'sd-2566}, {12'sd-1562, 11'sd708, 9'sd132}, {11'sd-648, 4'sd7, 11'sd922}},
{{12'sd-1436, 12'sd1220, 13'sd2564}, {12'sd1178, 9'sd161, 12'sd1680}, {11'sd-932, 13'sd2836, 11'sd-944}},
{{10'sd-339, 11'sd715, 12'sd1225}, {13'sd-2363, 13'sd-2971, 12'sd-1134}, {12'sd1347, 13'sd-2073, 13'sd-2136}},
{{12'sd1611, 11'sd-601, 13'sd2640}, {12'sd-1862, 10'sd-384, 9'sd-239}, {12'sd-1746, 11'sd1021, 12'sd1670}},
{{13'sd-2821, 12'sd1144, 11'sd979}, {12'sd1200, 12'sd1985, 13'sd2206}, {12'sd-1337, 10'sd-307, 13'sd3383}},
{{12'sd1192, 12'sd1507, 12'sd1660}, {13'sd2182, 10'sd-292, 10'sd-366}, {11'sd-919, 13'sd2433, 12'sd-2014}},
{{11'sd537, 10'sd397, 13'sd2275}, {12'sd1693, 12'sd1082, 11'sd-1002}, {12'sd1252, 12'sd1541, 13'sd-3172}},
{{12'sd1652, 12'sd-1025, 12'sd-1555}, {12'sd-1859, 8'sd96, 11'sd-1013}, {13'sd-2501, 12'sd-1846, 9'sd226}},
{{12'sd1328, 12'sd-1126, 12'sd1930}, {12'sd-1045, 12'sd-1083, 12'sd1493}, {11'sd-741, 12'sd1948, 12'sd1709}},
{{13'sd2915, 13'sd2231, 12'sd1131}, {12'sd1291, 9'sd-179, 12'sd1619}, {12'sd-1633, 11'sd-546, 13'sd-2965}},
{{13'sd-2411, 11'sd788, 11'sd-716}, {13'sd2888, 11'sd-582, 11'sd836}, {6'sd-28, 8'sd65, 10'sd-452}},
{{12'sd1468, 9'sd144, 10'sd483}, {12'sd1849, 13'sd-3001, 12'sd1885}, {10'sd360, 12'sd-1657, 13'sd-2882}},
{{12'sd1963, 13'sd2337, 12'sd-1215}, {10'sd-260, 11'sd-857, 12'sd1690}, {11'sd-601, 12'sd1593, 12'sd1620}},
{{7'sd-32, 13'sd-2659, 13'sd-2566}, {12'sd1081, 9'sd-137, 11'sd-995}, {11'sd-661, 7'sd-52, 12'sd-1928}},
{{10'sd304, 13'sd2076, 13'sd2400}, {13'sd2520, 13'sd2170, 11'sd524}, {13'sd2289, 9'sd152, 12'sd-1839}},
{{12'sd1118, 13'sd2329, 12'sd-1756}, {11'sd958, 13'sd2851, 12'sd1076}, {10'sd-396, 12'sd-1742, 12'sd-1048}},
{{10'sd451, 13'sd-3036, 13'sd2500}, {13'sd-2994, 12'sd1840, 11'sd-693}, {10'sd-432, 9'sd-250, 12'sd1276}},
{{12'sd-1375, 12'sd-1896, 12'sd1532}, {12'sd-1036, 12'sd-1864, 12'sd-1324}, {8'sd-106, 10'sd419, 11'sd-934}},
{{12'sd1603, 12'sd2015, 13'sd2490}, {13'sd2882, 12'sd-1985, 13'sd2709}, {13'sd2328, 12'sd-1099, 11'sd-944}},
{{6'sd-22, 12'sd-1212, 7'sd37}, {13'sd2699, 13'sd2297, 9'sd-162}, {10'sd-290, 12'sd2022, 13'sd2808}},
{{11'sd873, 12'sd1839, 12'sd-1407}, {10'sd327, 9'sd-143, 11'sd615}, {10'sd306, 9'sd232, 13'sd2209}},
{{9'sd-199, 13'sd-2182, 11'sd-590}, {9'sd155, 13'sd-2174, 12'sd1431}, {13'sd-2104, 10'sd-281, 12'sd-1576}},
{{11'sd-647, 12'sd1373, 11'sd-881}, {13'sd2317, 11'sd-524, 10'sd375}, {13'sd2510, 11'sd-781, 13'sd3383}},
{{12'sd1899, 9'sd241, 12'sd-1302}, {13'sd2546, 13'sd2551, 10'sd-382}, {12'sd-2031, 13'sd2306, 8'sd-92}},
{{13'sd-3578, 13'sd-2655, 10'sd-399}, {11'sd-919, 13'sd2277, 13'sd2536}, {13'sd-2157, 11'sd846, 9'sd-192}},
{{13'sd2197, 11'sd-856, 12'sd-1861}, {13'sd2593, 12'sd-1466, 13'sd-2886}, {10'sd-448, 12'sd1885, 12'sd1132}},
{{11'sd-632, 13'sd2398, 12'sd1247}, {13'sd-2319, 9'sd-150, 13'sd2513}, {11'sd934, 12'sd1559, 13'sd2083}},
{{13'sd2259, 13'sd-2736, 13'sd-2773}, {12'sd-1370, 11'sd740, 9'sd146}, {12'sd1874, 12'sd-1058, 12'sd-1910}},
{{12'sd-1314, 12'sd-1776, 9'sd-182}, {10'sd-450, 11'sd-885, 13'sd-2207}, {13'sd2102, 12'sd-1048, 12'sd1760}},
{{13'sd-2934, 13'sd-2946, 11'sd-759}, {11'sd776, 12'sd-1049, 12'sd1068}, {12'sd1452, 10'sd391, 13'sd2694}},
{{13'sd2124, 10'sd327, 11'sd-870}, {12'sd-1182, 13'sd2488, 12'sd1719}, {13'sd-3122, 12'sd-1230, 11'sd736}},
{{11'sd-561, 11'sd640, 12'sd1469}, {12'sd1537, 12'sd1028, 12'sd-1774}, {12'sd-1968, 13'sd-2182, 12'sd1669}},
{{12'sd1589, 12'sd-1681, 11'sd-955}, {12'sd-2004, 12'sd-1030, 13'sd2382}, {11'sd-612, 13'sd3232, 12'sd1804}},
{{13'sd-2143, 12'sd-1752, 11'sd-1016}, {13'sd-2691, 13'sd2115, 12'sd1809}, {10'sd-365, 12'sd1333, 10'sd460}},
{{13'sd2335, 12'sd2024, 12'sd-1270}, {12'sd-2043, 11'sd-906, 10'sd314}, {11'sd-841, 13'sd2956, 7'sd34}},
{{13'sd-2434, 12'sd-1855, 13'sd-2256}, {10'sd-402, 12'sd-2011, 12'sd-1495}, {13'sd-2125, 13'sd-2182, 11'sd-991}},
{{11'sd791, 12'sd1312, 12'sd-1089}, {11'sd-740, 13'sd3311, 6'sd-27}, {12'sd1864, 10'sd365, 12'sd-1169}},
{{12'sd1311, 12'sd1663, 12'sd-1573}, {12'sd1868, 12'sd1767, 9'sd211}, {11'sd695, 11'sd666, 13'sd-2785}},
{{11'sd681, 9'sd220, 10'sd-295}, {13'sd-2059, 11'sd-731, 13'sd-2598}, {7'sd41, 12'sd-1310, 12'sd1321}},
{{13'sd-2207, 12'sd-1737, 13'sd-2361}, {12'sd-1600, 12'sd-1596, 13'sd-2295}, {12'sd1227, 13'sd2510, 12'sd-1312}},
{{11'sd579, 11'sd630, 13'sd-3133}, {10'sd374, 12'sd-1066, 13'sd-3360}, {12'sd-1709, 11'sd-993, 13'sd-3302}},
{{13'sd3158, 12'sd-1638, 13'sd2077}, {11'sd906, 13'sd-2237, 4'sd7}, {13'sd2462, 8'sd105, 11'sd-723}},
{{13'sd-2463, 12'sd-1770, 12'sd1937}, {12'sd-1231, 13'sd2498, 13'sd2079}, {11'sd-676, 12'sd1169, 12'sd-1906}},
{{11'sd-848, 13'sd2936, 11'sd534}, {12'sd-1928, 11'sd-657, 12'sd1662}, {12'sd-1541, 12'sd-1242, 13'sd-2176}},
{{12'sd1617, 12'sd-1206, 13'sd-2339}, {12'sd-1689, 11'sd711, 13'sd-2190}, {12'sd-1610, 13'sd2579, 11'sd842}},
{{9'sd227, 12'sd-1540, 11'sd-631}, {13'sd-2322, 12'sd-1761, 12'sd-1572}, {11'sd795, 13'sd2842, 12'sd-1082}},
{{13'sd-3470, 11'sd-647, 13'sd-2327}, {13'sd-3202, 13'sd-2407, 11'sd885}, {11'sd634, 11'sd-955, 9'sd224}},
{{11'sd-775, 13'sd-2110, 13'sd2199}, {12'sd1777, 11'sd-781, 10'sd-436}, {11'sd-654, 12'sd-1504, 12'sd1729}},
{{11'sd542, 10'sd-308, 11'sd692}, {13'sd-2111, 11'sd-946, 13'sd2174}, {11'sd783, 6'sd-16, 13'sd-2815}},
{{11'sd859, 12'sd1662, 13'sd2429}, {13'sd2246, 13'sd2126, 13'sd2673}, {12'sd-1369, 11'sd961, 13'sd-2657}},
{{13'sd-2618, 10'sd283, 11'sd900}, {10'sd376, 13'sd2692, 11'sd818}, {12'sd1419, 12'sd-1776, 10'sd470}},
{{12'sd-1632, 12'sd2009, 10'sd349}, {6'sd22, 7'sd-37, 13'sd2443}, {13'sd2506, 11'sd-792, 9'sd191}},
{{13'sd2067, 11'sd598, 12'sd1907}, {12'sd1878, 12'sd1692, 11'sd722}, {10'sd366, 13'sd2145, 13'sd-2233}},
{{12'sd-1092, 13'sd-2845, 12'sd1369}, {13'sd2127, 13'sd-2583, 12'sd1866}, {12'sd-1761, 11'sd971, 11'sd1000}},
{{13'sd-3499, 13'sd-2623, 12'sd-1050}, {12'sd1955, 10'sd493, 12'sd-1289}, {13'sd-3305, 10'sd422, 10'sd-287}},
{{10'sd-479, 11'sd930, 11'sd917}, {13'sd2601, 13'sd-2345, 10'sd-302}, {11'sd-882, 12'sd1051, 13'sd-2174}}},
{
{{12'sd1177, 12'sd-1663, 13'sd2117}, {13'sd-2164, 11'sd-1001, 11'sd-843}, {10'sd-360, 11'sd607, 11'sd-531}},
{{11'sd808, 12'sd-1671, 10'sd424}, {13'sd2148, 13'sd2747, 8'sd-89}, {13'sd3357, 7'sd-62, 12'sd-1290}},
{{12'sd-1254, 10'sd259, 13'sd3078}, {10'sd353, 12'sd-1188, 11'sd693}, {13'sd-2781, 9'sd210, 12'sd-1818}},
{{7'sd50, 12'sd-1138, 13'sd3047}, {12'sd-1445, 9'sd-148, 10'sd408}, {11'sd-859, 11'sd-966, 13'sd2391}},
{{13'sd-3115, 9'sd-209, 12'sd1232}, {12'sd-1830, 12'sd1455, 13'sd-2558}, {11'sd915, 7'sd-59, 10'sd-339}},
{{13'sd-2364, 8'sd82, 12'sd-1750}, {9'sd249, 11'sd749, 13'sd2398}, {11'sd677, 12'sd-1281, 13'sd2091}},
{{10'sd395, 10'sd339, 12'sd-1358}, {11'sd625, 12'sd-1537, 9'sd-233}, {13'sd3110, 11'sd-602, 12'sd1535}},
{{13'sd2658, 12'sd1093, 12'sd1782}, {12'sd1970, 7'sd-45, 10'sd257}, {8'sd107, 12'sd1585, 10'sd-292}},
{{11'sd-966, 12'sd1581, 12'sd-1541}, {13'sd-3543, 12'sd-1363, 9'sd200}, {11'sd-678, 13'sd-2997, 11'sd-859}},
{{10'sd-324, 11'sd799, 8'sd-109}, {13'sd2654, 10'sd457, 11'sd591}, {12'sd1712, 13'sd2063, 12'sd1453}},
{{9'sd128, 13'sd2080, 12'sd1967}, {11'sd983, 7'sd33, 12'sd-1064}, {13'sd2123, 12'sd-1916, 6'sd-22}},
{{11'sd-560, 12'sd-1804, 11'sd-512}, {11'sd684, 12'sd1422, 11'sd-892}, {13'sd2067, 11'sd892, 10'sd344}},
{{12'sd1556, 12'sd-1792, 10'sd-426}, {12'sd1176, 11'sd-868, 12'sd-1419}, {12'sd1263, 13'sd-2476, 14'sd-4190}},
{{7'sd62, 13'sd2210, 9'sd221}, {13'sd2854, 12'sd1735, 12'sd-1418}, {6'sd-28, 11'sd-707, 13'sd2439}},
{{12'sd-1586, 6'sd-22, 12'sd1747}, {12'sd1619, 11'sd642, 14'sd4185}, {9'sd243, 13'sd2772, 13'sd3792}},
{{9'sd209, 10'sd-403, 13'sd2188}, {12'sd-1216, 13'sd2588, 11'sd787}, {11'sd747, 12'sd-1824, 11'sd-791}},
{{7'sd48, 12'sd-1744, 12'sd-1713}, {9'sd220, 12'sd1763, 13'sd-2586}, {12'sd1231, 11'sd996, 11'sd-539}},
{{14'sd-4676, 9'sd253, 13'sd-4060}, {13'sd-2864, 12'sd-1457, 13'sd-3330}, {13'sd-2330, 10'sd342, 13'sd-4004}},
{{13'sd2248, 12'sd1887, 12'sd-1148}, {11'sd583, 12'sd1914, 13'sd2139}, {12'sd-1154, 13'sd3539, 11'sd1012}},
{{12'sd1563, 12'sd-1407, 12'sd2026}, {13'sd-2278, 10'sd384, 12'sd1335}, {10'sd268, 13'sd-2659, 11'sd-832}},
{{11'sd551, 13'sd2134, 11'sd686}, {12'sd-1936, 12'sd1340, 11'sd827}, {13'sd-2772, 12'sd-1280, 11'sd843}},
{{13'sd2321, 12'sd-1883, 13'sd3434}, {12'sd1407, 10'sd281, 12'sd2010}, {11'sd705, 12'sd1116, 13'sd3141}},
{{10'sd-329, 13'sd2213, 13'sd2520}, {13'sd-2347, 13'sd3131, 11'sd786}, {13'sd-2353, 9'sd-246, 13'sd-3210}},
{{11'sd-852, 13'sd-2430, 12'sd1773}, {12'sd1348, 10'sd335, 12'sd1541}, {11'sd630, 3'sd-2, 10'sd273}},
{{12'sd-1685, 12'sd-1066, 11'sd-868}, {13'sd-2723, 13'sd-2241, 10'sd-336}, {12'sd1033, 12'sd1743, 11'sd522}},
{{11'sd683, 12'sd-1335, 12'sd-1351}, {12'sd1982, 11'sd977, 9'sd-145}, {13'sd-2129, 11'sd-667, 9'sd154}},
{{8'sd105, 11'sd-798, 10'sd311}, {11'sd931, 12'sd1666, 11'sd805}, {13'sd-2049, 7'sd63, 11'sd806}},
{{12'sd1507, 12'sd-1744, 12'sd1602}, {11'sd-739, 9'sd-151, 12'sd1857}, {13'sd2735, 13'sd2933, 12'sd1663}},
{{8'sd93, 12'sd-1116, 13'sd3050}, {12'sd-1566, 9'sd-195, 10'sd-274}, {10'sd-502, 9'sd236, 12'sd1542}},
{{11'sd-642, 10'sd258, 12'sd1441}, {11'sd-579, 13'sd2267, 12'sd1372}, {12'sd1844, 5'sd12, 7'sd-48}},
{{12'sd-1268, 12'sd-1247, 12'sd-1573}, {11'sd-628, 10'sd411, 12'sd-1392}, {13'sd3293, 12'sd1272, 9'sd195}},
{{12'sd-1238, 9'sd180, 12'sd-1531}, {12'sd1351, 11'sd-860, 13'sd-2622}, {9'sd144, 12'sd-1773, 13'sd-2862}},
{{9'sd212, 12'sd-1700, 13'sd-2785}, {12'sd1843, 9'sd249, 11'sd-922}, {11'sd911, 7'sd62, 14'sd-5048}},
{{11'sd-730, 11'sd804, 13'sd2139}, {13'sd2819, 10'sd414, 13'sd2267}, {11'sd571, 13'sd2685, 11'sd595}},
{{12'sd1804, 1'sd0, 12'sd1326}, {13'sd2665, 12'sd-1949, 12'sd1528}, {11'sd841, 12'sd1331, 10'sd264}},
{{9'sd-187, 11'sd833, 13'sd2339}, {12'sd-1686, 11'sd688, 12'sd1953}, {10'sd343, 10'sd354, 11'sd-600}},
{{11'sd924, 6'sd25, 12'sd1936}, {10'sd-478, 10'sd465, 11'sd-956}, {12'sd1723, 12'sd1755, 13'sd2073}},
{{12'sd1696, 12'sd-1788, 13'sd2237}, {12'sd1357, 13'sd2076, 12'sd-1451}, {12'sd-1362, 12'sd1954, 12'sd1586}},
{{12'sd-1276, 12'sd-1816, 13'sd2916}, {12'sd-1679, 13'sd2155, 7'sd-40}, {13'sd-2421, 12'sd1140, 11'sd-599}},
{{3'sd-2, 11'sd-813, 13'sd2317}, {10'sd268, 12'sd1585, 12'sd-1942}, {11'sd-989, 12'sd1247, 12'sd-1646}},
{{11'sd-839, 10'sd-393, 9'sd-191}, {13'sd-2828, 13'sd2617, 12'sd-1316}, {12'sd-1206, 13'sd-2494, 12'sd-1692}},
{{11'sd556, 10'sd503, 12'sd-1264}, {10'sd-274, 12'sd-1387, 12'sd-1460}, {13'sd-2319, 13'sd-2201, 9'sd-148}},
{{12'sd-1692, 11'sd881, 10'sd-322}, {13'sd-2284, 10'sd-317, 12'sd-1134}, {13'sd-2400, 11'sd-544, 13'sd-3122}},
{{12'sd-1505, 13'sd-2746, 11'sd674}, {10'sd-368, 12'sd-1927, 12'sd1774}, {13'sd-2537, 12'sd1646, 10'sd-265}},
{{13'sd-2591, 8'sd87, 12'sd-1519}, {12'sd-1790, 10'sd-276, 12'sd-2032}, {12'sd-2016, 12'sd-1934, 12'sd1365}},
{{12'sd1126, 11'sd945, 9'sd179}, {13'sd-2665, 8'sd-93, 13'sd-2265}, {11'sd-559, 7'sd-48, 12'sd1353}},
{{12'sd1339, 12'sd-1285, 13'sd2544}, {10'sd-345, 10'sd-366, 12'sd1300}, {13'sd-2976, 12'sd-1735, 12'sd1637}},
{{11'sd822, 13'sd-2335, 11'sd-663}, {11'sd1012, 12'sd-2035, 11'sd-853}, {12'sd1489, 11'sd856, 13'sd2204}},
{{12'sd1181, 12'sd1340, 10'sd-414}, {10'sd434, 13'sd3893, 12'sd-2046}, {13'sd2874, 11'sd778, 13'sd-2848}},
{{12'sd-1392, 12'sd1565, 12'sd-2032}, {13'sd-3369, 12'sd-1026, 7'sd62}, {11'sd-1019, 13'sd3179, 10'sd-342}},
{{13'sd3466, 13'sd-2227, 10'sd-297}, {13'sd2262, 12'sd1537, 13'sd2208}, {14'sd-4680, 13'sd-2996, 12'sd-1369}},
{{13'sd-2254, 11'sd975, 10'sd-465}, {11'sd-1016, 13'sd-2638, 12'sd-1822}, {12'sd1250, 13'sd-3175, 12'sd-1070}},
{{9'sd241, 12'sd1699, 13'sd-2291}, {11'sd-962, 11'sd839, 12'sd-1532}, {12'sd1721, 10'sd285, 11'sd-599}},
{{13'sd-3008, 10'sd-266, 10'sd-435}, {12'sd-1395, 12'sd-1423, 12'sd1084}, {10'sd-459, 10'sd363, 13'sd2102}},
{{12'sd-1729, 12'sd-1404, 12'sd-1372}, {12'sd-1425, 13'sd-2085, 11'sd-580}, {7'sd38, 13'sd-3790, 14'sd-4234}},
{{12'sd1110, 12'sd-1309, 11'sd907}, {13'sd2325, 13'sd2398, 13'sd2212}, {11'sd-682, 11'sd985, 9'sd-246}},
{{12'sd1335, 13'sd2679, 13'sd3384}, {11'sd779, 10'sd348, 11'sd988}, {9'sd-133, 13'sd3263, 11'sd687}},
{{10'sd-418, 12'sd1781, 9'sd236}, {11'sd574, 13'sd2164, 12'sd1621}, {14'sd4173, 13'sd2884, 13'sd3256}},
{{13'sd3497, 13'sd-2081, 11'sd-562}, {13'sd2595, 12'sd-1557, 12'sd-1834}, {12'sd1237, 12'sd-1376, 11'sd817}},
{{11'sd-677, 12'sd1262, 13'sd2593}, {13'sd2447, 11'sd998, 11'sd-867}, {12'sd1719, 13'sd-2122, 11'sd-766}},
{{13'sd-2919, 12'sd1615, 11'sd583}, {13'sd-2295, 11'sd929, 9'sd-221}, {13'sd-2283, 12'sd1930, 13'sd2480}},
{{11'sd549, 12'sd-2009, 11'sd-530}, {13'sd2565, 13'sd2735, 13'sd-2264}, {13'sd3679, 13'sd3776, 13'sd-2976}},
{{6'sd-21, 10'sd484, 13'sd3114}, {12'sd-1356, 12'sd-1459, 11'sd653}, {11'sd684, 10'sd-460, 12'sd1933}},
{{11'sd769, 11'sd-854, 12'sd-1838}, {13'sd-2287, 13'sd-2131, 10'sd492}, {11'sd-615, 13'sd2503, 13'sd-2493}}},
{
{{11'sd-762, 9'sd170, 12'sd1089}, {13'sd-2082, 13'sd-2358, 11'sd-837}, {12'sd-1755, 13'sd-2096, 12'sd1745}},
{{12'sd-1547, 11'sd-516, 12'sd1262}, {12'sd1092, 12'sd1304, 9'sd-243}, {12'sd1604, 13'sd-2725, 12'sd-1948}},
{{12'sd-1595, 10'sd390, 13'sd3062}, {12'sd-1276, 9'sd-206, 12'sd-1583}, {14'sd-4249, 12'sd-1074, 12'sd-1883}},
{{8'sd118, 8'sd-126, 13'sd-2911}, {8'sd-118, 13'sd-3537, 13'sd-3027}, {13'sd2156, 13'sd-3416, 12'sd1199}},
{{13'sd2286, 12'sd-1607, 12'sd2044}, {12'sd1426, 13'sd2666, 12'sd1283}, {12'sd1490, 13'sd2239, 12'sd1920}},
{{12'sd-1114, 12'sd-1770, 13'sd2413}, {12'sd1157, 12'sd1912, 12'sd-1133}, {13'sd-2303, 12'sd-1817, 13'sd2525}},
{{10'sd-275, 13'sd-3204, 12'sd1713}, {12'sd-1289, 12'sd-1898, 13'sd-2247}, {13'sd3623, 10'sd-308, 8'sd-109}},
{{14'sd-4302, 13'sd-2580, 14'sd-4831}, {12'sd-1200, 11'sd873, 13'sd-2965}, {11'sd-643, 12'sd1566, 8'sd-116}},
{{8'sd-118, 13'sd-2458, 12'sd1052}, {13'sd2296, 11'sd-941, 13'sd-2306}, {13'sd2638, 13'sd-3485, 10'sd344}},
{{12'sd1457, 7'sd-54, 8'sd66}, {12'sd-1863, 12'sd1421, 12'sd1987}, {13'sd2417, 10'sd-328, 10'sd289}},
{{13'sd2095, 11'sd709, 13'sd2184}, {11'sd-749, 9'sd240, 13'sd2715}, {13'sd2552, 12'sd-1839, 12'sd-1651}},
{{13'sd-2130, 11'sd560, 11'sd731}, {9'sd225, 11'sd516, 11'sd-801}, {12'sd1058, 11'sd-594, 6'sd-24}},
{{12'sd-1565, 13'sd-2783, 12'sd1292}, {11'sd-939, 13'sd-2868, 13'sd-2939}, {12'sd1636, 5'sd-14, 9'sd-214}},
{{12'sd-1044, 6'sd-26, 12'sd-1287}, {13'sd-2378, 12'sd-1987, 11'sd-964}, {9'sd153, 12'sd-1148, 12'sd1850}},
{{10'sd-310, 11'sd910, 12'sd1359}, {13'sd-2546, 13'sd2164, 12'sd-1920}, {12'sd1466, 13'sd-2779, 12'sd-1315}},
{{13'sd2516, 13'sd2758, 12'sd1937}, {10'sd283, 12'sd1335, 12'sd-1756}, {12'sd1495, 12'sd-1259, 12'sd1135}},
{{11'sd788, 13'sd-2088, 10'sd429}, {12'sd1956, 11'sd-709, 10'sd-310}, {11'sd677, 12'sd1123, 13'sd-2267}},
{{11'sd685, 12'sd1250, 13'sd-2766}, {13'sd2841, 13'sd-2298, 13'sd-3292}, {11'sd-613, 13'sd-2490, 13'sd-3397}},
{{13'sd-2349, 11'sd763, 11'sd-803}, {10'sd-482, 13'sd2471, 13'sd-2048}, {11'sd-965, 12'sd1268, 13'sd-3064}},
{{10'sd299, 12'sd1256, 12'sd-1689}, {11'sd-725, 11'sd982, 12'sd1334}, {12'sd-1144, 12'sd1225, 12'sd1362}},
{{11'sd-680, 11'sd-754, 10'sd-323}, {11'sd-670, 10'sd-282, 12'sd1361}, {10'sd442, 13'sd2684, 13'sd3027}},
{{12'sd1271, 9'sd198, 12'sd1160}, {8'sd76, 13'sd-2929, 11'sd-936}, {12'sd1208, 10'sd-477, 12'sd-1502}},
{{7'sd35, 11'sd-658, 13'sd-2269}, {13'sd-2465, 12'sd1161, 10'sd487}, {11'sd897, 10'sd-444, 12'sd1283}},
{{12'sd1769, 12'sd-1277, 11'sd-749}, {9'sd-177, 12'sd-1842, 12'sd-1519}, {12'sd1699, 8'sd-65, 11'sd617}},
{{12'sd-1937, 12'sd-1683, 13'sd2247}, {13'sd2577, 11'sd1001, 11'sd-869}, {11'sd890, 10'sd-508, 12'sd-1794}},
{{12'sd-1520, 13'sd-2144, 12'sd-1900}, {12'sd1683, 9'sd171, 11'sd1003}, {11'sd-954, 12'sd1503, 13'sd2952}},
{{9'sd-224, 12'sd1710, 12'sd1907}, {12'sd1098, 11'sd-757, 3'sd3}, {13'sd-2159, 11'sd546, 11'sd855}},
{{12'sd1281, 12'sd-1575, 13'sd-2089}, {12'sd1651, 10'sd388, 11'sd976}, {12'sd-1849, 10'sd323, 12'sd-1220}},
{{12'sd-1135, 11'sd-697, 13'sd3577}, {13'sd-2218, 12'sd-1171, 13'sd3325}, {12'sd-1084, 10'sd-479, 11'sd-572}},
{{13'sd-2868, 12'sd1427, 12'sd-1297}, {11'sd957, 12'sd1131, 9'sd157}, {13'sd-2404, 11'sd658, 12'sd-1309}},
{{11'sd974, 11'sd905, 11'sd-647}, {12'sd1830, 13'sd2715, 13'sd2337}, {9'sd-163, 13'sd3911, 12'sd-1246}},
{{11'sd-652, 12'sd1878, 13'sd2447}, {9'sd-190, 13'sd2335, 11'sd591}, {7'sd52, 13'sd-2629, 13'sd-2700}},
{{14'sd-4153, 12'sd-1329, 13'sd-2700}, {11'sd638, 13'sd2592, 12'sd1077}, {11'sd-681, 13'sd-2059, 13'sd3289}},
{{11'sd-1016, 11'sd-937, 13'sd2465}, {12'sd1175, 10'sd324, 12'sd1701}, {10'sd-403, 13'sd2699, 13'sd-2647}},
{{12'sd-1362, 13'sd-2601, 13'sd2111}, {13'sd-2890, 13'sd-2462, 10'sd421}, {12'sd1414, 12'sd-1107, 12'sd-1222}},
{{12'sd-1639, 12'sd1576, 10'sd-484}, {12'sd-1362, 13'sd-2567, 12'sd-1125}, {13'sd-2415, 12'sd1242, 13'sd-2058}},
{{7'sd-37, 13'sd2517, 12'sd-1846}, {9'sd186, 12'sd-1291, 12'sd2003}, {12'sd-1660, 12'sd-1205, 12'sd-1403}},
{{12'sd-1670, 12'sd1507, 12'sd-1475}, {12'sd1707, 12'sd1609, 10'sd-310}, {11'sd571, 12'sd1674, 12'sd-1106}},
{{11'sd1009, 8'sd79, 8'sd80}, {12'sd-2016, 13'sd-2129, 12'sd1502}, {11'sd-697, 12'sd1453, 12'sd1986}},
{{7'sd53, 11'sd1001, 12'sd-1663}, {12'sd1505, 11'sd597, 12'sd1296}, {10'sd441, 8'sd-117, 12'sd-1210}},
{{11'sd602, 11'sd-551, 7'sd40}, {12'sd-1488, 12'sd1361, 5'sd-12}, {9'sd-206, 13'sd3204, 12'sd1942}},
{{11'sd-800, 12'sd1327, 13'sd2999}, {13'sd-2781, 10'sd-302, 11'sd732}, {10'sd496, 12'sd-1800, 11'sd-982}},
{{12'sd1656, 11'sd-855, 12'sd-1116}, {11'sd666, 10'sd-485, 13'sd2730}, {9'sd-223, 12'sd1411, 12'sd-1167}},
{{13'sd-2657, 13'sd-2766, 12'sd-1186}, {12'sd1065, 12'sd1898, 10'sd-350}, {13'sd2392, 13'sd2513, 13'sd-2058}},
{{13'sd-2194, 13'sd-2294, 11'sd-904}, {11'sd526, 11'sd723, 10'sd-293}, {13'sd-2902, 11'sd-807, 13'sd2252}},
{{13'sd-2184, 10'sd342, 12'sd-1145}, {5'sd14, 9'sd134, 12'sd1415}, {11'sd-519, 12'sd1313, 12'sd-1093}},
{{12'sd1219, 11'sd973, 13'sd2390}, {13'sd-3156, 8'sd90, 9'sd250}, {11'sd-521, 11'sd719, 11'sd-590}},
{{12'sd-1336, 11'sd-545, 8'sd-82}, {11'sd-773, 11'sd-880, 12'sd1689}, {11'sd-819, 12'sd-1973, 9'sd-141}},
{{12'sd1876, 12'sd-1572, 12'sd-1209}, {12'sd-1397, 13'sd2296, 13'sd-2189}, {12'sd1798, 11'sd736, 11'sd925}},
{{12'sd-1588, 11'sd560, 13'sd-3225}, {13'sd-2632, 13'sd2574, 11'sd-916}, {13'sd-2606, 12'sd1069, 9'sd-148}},
{{13'sd-2735, 13'sd2459, 13'sd2294}, {9'sd155, 12'sd1243, 13'sd3023}, {13'sd-3267, 12'sd1433, 12'sd1952}},
{{11'sd-541, 12'sd-1376, 13'sd-2229}, {12'sd-1254, 12'sd-1068, 10'sd-467}, {13'sd-2748, 12'sd1818, 12'sd1976}},
{{13'sd-2232, 12'sd1196, 13'sd2860}, {11'sd-579, 13'sd-2400, 11'sd572}, {10'sd-281, 8'sd-125, 11'sd-958}},
{{13'sd-2287, 10'sd411, 10'sd511}, {11'sd722, 11'sd-844, 12'sd-1064}, {13'sd-2703, 13'sd2340, 12'sd1301}},
{{12'sd1343, 7'sd-35, 12'sd1802}, {11'sd605, 13'sd2907, 12'sd-1203}, {11'sd-716, 12'sd1077, 13'sd-2237}},
{{13'sd2184, 9'sd-233, 7'sd44}, {11'sd822, 13'sd-2179, 13'sd-2212}, {12'sd1453, 10'sd452, 13'sd-2299}},
{{10'sd-349, 12'sd1254, 11'sd852}, {13'sd-2048, 11'sd713, 11'sd873}, {12'sd1620, 11'sd-954, 10'sd-422}},
{{12'sd1408, 13'sd2687, 12'sd-1625}, {6'sd28, 12'sd-1679, 11'sd-863}, {12'sd1237, 12'sd-1979, 11'sd602}},
{{13'sd-2059, 8'sd-64, 13'sd-2104}, {12'sd-1219, 12'sd-1517, 13'sd2131}, {13'sd2856, 7'sd40, 13'sd2345}},
{{13'sd3753, 13'sd-2139, 11'sd902}, {13'sd2446, 12'sd-1495, 10'sd459}, {8'sd-127, 12'sd-1189, 9'sd-176}},
{{11'sd1013, 12'sd1486, 12'sd1148}, {10'sd-340, 11'sd-690, 12'sd-1392}, {10'sd357, 12'sd1170, 12'sd1702}},
{{13'sd-3128, 8'sd-108, 12'sd1681}, {12'sd1596, 12'sd-1036, 11'sd885}, {12'sd1163, 12'sd1814, 12'sd1422}},
{{11'sd-791, 10'sd-345, 7'sd61}, {12'sd1929, 13'sd3105, 11'sd-798}, {12'sd1665, 13'sd2793, 12'sd-1208}},
{{11'sd958, 12'sd-1418, 8'sd76}, {11'sd897, 12'sd-1808, 13'sd-2937}, {12'sd-1582, 10'sd386, 12'sd-1486}}},
{
{{13'sd-2769, 12'sd1257, 13'sd2186}, {11'sd-794, 10'sd-469, 13'sd2173}, {12'sd-1432, 13'sd-2119, 12'sd1932}},
{{13'sd-2428, 10'sd-339, 13'sd-2505}, {13'sd-2245, 13'sd-2382, 13'sd-2675}, {13'sd-2629, 13'sd-2119, 12'sd1677}},
{{13'sd3120, 12'sd1040, 12'sd1474}, {12'sd-1881, 10'sd354, 12'sd-1653}, {13'sd-2280, 12'sd1172, 12'sd1245}},
{{13'sd-2666, 12'sd1247, 11'sd776}, {11'sd770, 11'sd856, 13'sd-2761}, {11'sd900, 13'sd-2266, 10'sd302}},
{{12'sd2013, 13'sd-2161, 12'sd1397}, {12'sd1909, 12'sd1702, 13'sd2319}, {11'sd589, 12'sd-1152, 13'sd2309}},
{{12'sd-1663, 10'sd-384, 12'sd-1306}, {12'sd-1042, 12'sd1193, 12'sd1810}, {13'sd-2134, 13'sd2354, 13'sd-2760}},
{{13'sd3065, 13'sd-2713, 10'sd-447}, {11'sd1008, 12'sd-1173, 12'sd-1592}, {12'sd-1526, 10'sd507, 13'sd-2933}},
{{11'sd-1014, 12'sd-1562, 12'sd-1330}, {12'sd1998, 12'sd-1985, 12'sd-1289}, {10'sd-432, 10'sd369, 13'sd-2919}},
{{11'sd761, 10'sd-269, 11'sd-993}, {11'sd564, 12'sd-1964, 10'sd-371}, {13'sd2497, 12'sd2027, 13'sd-2617}},
{{13'sd-2187, 12'sd1852, 10'sd-278}, {10'sd-445, 12'sd1940, 12'sd1424}, {7'sd53, 13'sd-2108, 12'sd1488}},
{{12'sd-1065, 13'sd-2144, 12'sd1444}, {11'sd-998, 13'sd3252, 12'sd1349}, {11'sd563, 11'sd-557, 10'sd-458}},
{{12'sd-1691, 12'sd-1148, 10'sd387}, {12'sd-1103, 12'sd-1492, 10'sd-308}, {10'sd-325, 11'sd965, 13'sd-2694}},
{{12'sd-1186, 13'sd2625, 9'sd198}, {12'sd1190, 11'sd-1003, 10'sd351}, {13'sd-2737, 11'sd564, 12'sd-1686}},
{{10'sd441, 13'sd2186, 12'sd-1708}, {11'sd810, 11'sd862, 13'sd-2159}, {9'sd233, 11'sd-679, 10'sd-399}},
{{12'sd-1312, 13'sd2483, 11'sd613}, {13'sd2524, 12'sd1043, 12'sd1872}, {13'sd2605, 12'sd-1085, 12'sd-1872}},
{{13'sd-2246, 12'sd-1538, 12'sd2026}, {9'sd161, 13'sd2268, 12'sd1819}, {12'sd-1258, 11'sd575, 13'sd-2175}},
{{11'sd-830, 13'sd-2241, 13'sd2048}, {13'sd-2273, 12'sd-1968, 6'sd-17}, {10'sd-362, 10'sd356, 10'sd-360}},
{{10'sd-400, 6'sd-28, 11'sd631}, {10'sd417, 13'sd3526, 11'sd-907}, {11'sd-597, 12'sd1918, 13'sd3031}},
{{6'sd28, 12'sd-1981, 13'sd2574}, {10'sd388, 11'sd-789, 12'sd1580}, {12'sd-1329, 12'sd1374, 12'sd2036}},
{{12'sd-1253, 12'sd-1206, 13'sd-2157}, {12'sd1884, 11'sd-573, 10'sd357}, {12'sd-1561, 10'sd-312, 12'sd1175}},
{{11'sd-608, 13'sd2917, 13'sd-2287}, {12'sd1731, 12'sd1858, 10'sd287}, {12'sd-1310, 11'sd-632, 9'sd-195}},
{{13'sd-2688, 9'sd-252, 11'sd998}, {13'sd2713, 9'sd151, 12'sd-1102}, {13'sd-2790, 11'sd623, 12'sd1182}},
{{12'sd1427, 12'sd-1171, 11'sd945}, {12'sd1662, 7'sd-47, 10'sd-298}, {12'sd-2004, 12'sd1852, 9'sd164}},
{{10'sd473, 13'sd-2695, 13'sd-2776}, {9'sd-241, 13'sd-2347, 13'sd-2134}, {13'sd-2887, 12'sd1993, 13'sd-2590}},
{{12'sd1374, 10'sd324, 13'sd-2392}, {10'sd443, 12'sd1217, 13'sd2810}, {12'sd1543, 10'sd-428, 12'sd-1906}},
{{9'sd225, 12'sd-1606, 12'sd-1636}, {13'sd2255, 9'sd-153, 13'sd2506}, {11'sd-788, 11'sd-516, 13'sd2974}},
{{11'sd576, 12'sd2034, 9'sd194}, {8'sd-123, 12'sd1538, 13'sd-2262}, {11'sd614, 11'sd966, 12'sd-1066}},
{{11'sd640, 12'sd1854, 13'sd-2588}, {12'sd-1425, 10'sd257, 13'sd-2754}, {11'sd-997, 12'sd-1941, 13'sd2125}},
{{13'sd2073, 13'sd-2291, 11'sd-1004}, {13'sd-2054, 13'sd-2569, 11'sd925}, {10'sd-281, 13'sd2319, 12'sd1899}},
{{11'sd541, 12'sd1718, 13'sd2375}, {12'sd1629, 12'sd-1464, 13'sd-2492}, {12'sd1961, 7'sd54, 10'sd311}},
{{10'sd-406, 11'sd-823, 12'sd1536}, {12'sd-1242, 12'sd1178, 14'sd4240}, {14'sd-4549, 13'sd-2113, 12'sd-1304}},
{{13'sd-2203, 12'sd1234, 12'sd1881}, {13'sd-2614, 12'sd-1857, 9'sd223}, {12'sd1650, 12'sd1632, 13'sd-2056}},
{{11'sd-925, 9'sd240, 12'sd1576}, {12'sd-1810, 11'sd-537, 13'sd-2111}, {8'sd70, 13'sd2049, 10'sd-304}},
{{11'sd-590, 12'sd1055, 11'sd-561}, {10'sd484, 8'sd-89, 12'sd2019}, {12'sd1790, 10'sd-458, 13'sd-2244}},
{{12'sd-1873, 9'sd-178, 13'sd2436}, {12'sd1143, 12'sd-1440, 11'sd-716}, {13'sd2707, 12'sd-1954, 11'sd857}},
{{12'sd1463, 10'sd-420, 11'sd-890}, {12'sd-1522, 12'sd1829, 7'sd63}, {12'sd1801, 12'sd-1418, 12'sd1370}},
{{12'sd1068, 12'sd-1375, 12'sd-1761}, {11'sd-612, 12'sd-1273, 9'sd194}, {12'sd-1579, 13'sd2280, 13'sd-2758}},
{{13'sd2075, 11'sd-878, 11'sd810}, {10'sd295, 11'sd707, 13'sd2376}, {11'sd-538, 3'sd-3, 12'sd-1122}},
{{12'sd1776, 12'sd1221, 13'sd2532}, {13'sd-2557, 13'sd2078, 12'sd1199}, {9'sd-246, 11'sd615, 13'sd-2295}},
{{13'sd-2786, 10'sd264, 11'sd-659}, {13'sd-2667, 12'sd1979, 11'sd843}, {11'sd837, 8'sd100, 12'sd-1153}},
{{13'sd2694, 11'sd1003, 13'sd2259}, {13'sd2318, 12'sd-1272, 11'sd820}, {11'sd-789, 11'sd875, 12'sd1108}},
{{6'sd23, 12'sd-1583, 8'sd-81}, {10'sd373, 12'sd-1309, 13'sd-2681}, {13'sd2601, 9'sd-251, 13'sd2694}},
{{11'sd-1006, 8'sd86, 13'sd2608}, {9'sd130, 9'sd-213, 12'sd1400}, {10'sd-491, 11'sd-593, 12'sd-1121}},
{{12'sd-1782, 12'sd2003, 10'sd-450}, {13'sd2251, 11'sd597, 13'sd3017}, {13'sd3042, 13'sd2739, 12'sd-1486}},
{{11'sd-853, 12'sd1581, 12'sd-1929}, {13'sd2967, 12'sd-1946, 12'sd1307}, {12'sd1764, 12'sd-1252, 13'sd-2427}},
{{13'sd2891, 11'sd807, 12'sd1446}, {13'sd-2103, 11'sd-919, 13'sd2864}, {13'sd2418, 12'sd1530, 12'sd1215}},
{{12'sd1986, 13'sd-2248, 13'sd2742}, {10'sd305, 13'sd3190, 10'sd332}, {12'sd-1940, 13'sd2703, 9'sd-139}},
{{9'sd-164, 12'sd1033, 11'sd922}, {12'sd-1344, 13'sd-3419, 13'sd-2668}, {12'sd1719, 12'sd-1282, 13'sd-3566}},
{{3'sd-2, 13'sd3000, 13'sd2226}, {12'sd1669, 11'sd955, 12'sd1551}, {11'sd915, 12'sd-1675, 13'sd-2390}},
{{12'sd-1568, 10'sd453, 13'sd2400}, {12'sd1365, 6'sd20, 12'sd1026}, {11'sd-690, 13'sd2663, 12'sd-1993}},
{{11'sd-576, 13'sd2113, 13'sd2194}, {12'sd1755, 13'sd-2891, 11'sd-777}, {12'sd1409, 13'sd-2357, 8'sd-88}},
{{13'sd-2468, 11'sd-589, 12'sd-1940}, {12'sd1783, 13'sd-2799, 10'sd-365}, {13'sd2291, 10'sd-483, 12'sd-1608}},
{{11'sd-897, 12'sd-1751, 12'sd-1488}, {11'sd-735, 12'sd-1141, 12'sd-1782}, {13'sd2318, 12'sd1175, 8'sd72}},
{{13'sd-2786, 11'sd-1008, 13'sd2425}, {13'sd-2392, 12'sd-1840, 13'sd-2335}, {13'sd2271, 13'sd2168, 11'sd724}},
{{12'sd-1302, 11'sd961, 8'sd-85}, {11'sd1010, 12'sd-1546, 12'sd1224}, {13'sd-2409, 13'sd-2126, 10'sd458}},
{{7'sd-39, 13'sd-2333, 12'sd1295}, {13'sd2326, 13'sd-2152, 9'sd199}, {13'sd2758, 10'sd-312, 13'sd2843}},
{{11'sd542, 12'sd-1783, 11'sd597}, {9'sd-161, 13'sd2207, 12'sd-1160}, {10'sd-461, 11'sd834, 12'sd-1624}},
{{11'sd931, 12'sd2003, 11'sd722}, {11'sd818, 13'sd2844, 11'sd-985}, {12'sd1689, 12'sd-2035, 12'sd1065}},
{{12'sd-1478, 12'sd-1025, 12'sd1319}, {11'sd830, 11'sd553, 13'sd-2676}, {11'sd626, 13'sd-2698, 13'sd2712}},
{{13'sd2754, 12'sd-1187, 12'sd-1037}, {12'sd-1528, 12'sd1758, 10'sd-446}, {13'sd-2236, 12'sd1516, 12'sd-2047}},
{{9'sd-192, 11'sd-680, 11'sd-914}, {10'sd-319, 10'sd490, 13'sd2432}, {11'sd531, 12'sd-1412, 13'sd2336}},
{{12'sd1478, 12'sd-1921, 11'sd792}, {12'sd-2044, 13'sd2181, 13'sd2532}, {10'sd-334, 11'sd735, 12'sd-1926}},
{{11'sd884, 11'sd-634, 12'sd-1279}, {11'sd-689, 11'sd-707, 8'sd-83}, {13'sd-2233, 12'sd1359, 12'sd-1477}},
{{11'sd-732, 12'sd-1596, 9'sd249}, {11'sd598, 11'sd-582, 12'sd1246}, {13'sd-2113, 10'sd266, 13'sd-2318}}},
{
{{11'sd-582, 13'sd2533, 11'sd573}, {12'sd-1335, 13'sd-2977, 12'sd-1803}, {13'sd2375, 9'sd-133, 13'sd2696}},
{{12'sd-1493, 10'sd-476, 11'sd802}, {13'sd-2090, 11'sd798, 10'sd-420}, {12'sd-1333, 12'sd-1044, 12'sd1669}},
{{13'sd2434, 10'sd-440, 10'sd324}, {10'sd-478, 10'sd-509, 13'sd-2424}, {12'sd1578, 12'sd1954, 14'sd5315}},
{{12'sd-1386, 11'sd618, 13'sd-2952}, {5'sd-15, 13'sd-2059, 12'sd-1054}, {13'sd-3254, 14'sd-4320, 14'sd-5282}},
{{13'sd2614, 13'sd2853, 10'sd375}, {11'sd-911, 10'sd-423, 12'sd-1533}, {13'sd-2508, 12'sd-1693, 12'sd-1349}},
{{13'sd2879, 12'sd-1416, 12'sd1782}, {13'sd-2216, 11'sd959, 11'sd575}, {12'sd-1383, 12'sd1095, 13'sd2274}},
{{11'sd773, 13'sd-2527, 12'sd1949}, {12'sd-1803, 13'sd-2160, 12'sd-1668}, {12'sd1621, 13'sd3359, 12'sd-1174}},
{{12'sd1224, 12'sd1938, 11'sd623}, {13'sd-2954, 9'sd174, 12'sd-1972}, {12'sd-1277, 11'sd-785, 11'sd562}},
{{13'sd3362, 10'sd511, 9'sd-135}, {11'sd-758, 8'sd-100, 12'sd1591}, {13'sd2051, 12'sd-1598, 13'sd-2428}},
{{12'sd1508, 10'sd-385, 13'sd-2542}, {12'sd-1352, 13'sd-2067, 10'sd-441}, {13'sd3084, 13'sd-2074, 12'sd-1214}},
{{12'sd-1177, 10'sd-374, 12'sd-1125}, {11'sd-639, 13'sd2076, 12'sd1711}, {12'sd-1797, 11'sd-779, 4'sd-6}},
{{12'sd1845, 12'sd1720, 13'sd-2266}, {12'sd-1521, 12'sd-1640, 11'sd-597}, {12'sd1508, 12'sd1693, 13'sd3173}},
{{12'sd-1497, 2'sd-1, 13'sd-2257}, {13'sd3157, 10'sd-432, 11'sd604}, {11'sd615, 10'sd256, 12'sd1975}},
{{10'sd-398, 12'sd1936, 13'sd-2622}, {9'sd-244, 13'sd2278, 12'sd-1721}, {13'sd2410, 11'sd621, 10'sd389}},
{{11'sd602, 12'sd-1836, 12'sd-1210}, {11'sd1016, 13'sd-2858, 10'sd-431}, {13'sd-2554, 12'sd1475, 13'sd-3430}},
{{13'sd-2472, 11'sd-851, 12'sd-1104}, {8'sd-105, 12'sd-1943, 11'sd-709}, {12'sd1419, 13'sd2528, 13'sd3097}},
{{12'sd-2019, 13'sd-2266, 12'sd-1630}, {13'sd-2460, 12'sd-1576, 12'sd-1077}, {13'sd2114, 9'sd203, 12'sd1871}},
{{11'sd-862, 11'sd937, 12'sd2027}, {13'sd2877, 12'sd-1771, 11'sd-931}, {14'sd4966, 12'sd-1843, 10'sd-398}},
{{12'sd1968, 13'sd-3820, 11'sd-983}, {9'sd-245, 13'sd-3022, 11'sd783}, {9'sd-149, 12'sd-1221, 11'sd-567}},
{{10'sd472, 8'sd-68, 10'sd-451}, {11'sd-982, 3'sd3, 12'sd-1174}, {12'sd-1201, 12'sd1768, 13'sd2802}},
{{13'sd2160, 10'sd511, 13'sd-3830}, {12'sd-1404, 12'sd1293, 13'sd-2725}, {13'sd-2594, 13'sd-2649, 12'sd-1416}},
{{12'sd1599, 12'sd-1600, 9'sd239}, {12'sd1524, 9'sd164, 10'sd433}, {11'sd652, 13'sd3394, 12'sd1656}},
{{13'sd2178, 12'sd1174, 11'sd-808}, {11'sd-963, 12'sd1396, 13'sd-2409}, {9'sd-178, 11'sd1018, 10'sd-326}},
{{7'sd-52, 13'sd-2072, 13'sd2068}, {11'sd-596, 11'sd780, 13'sd-2394}, {13'sd-2783, 5'sd-11, 12'sd-1426}},
{{13'sd-2940, 11'sd-684, 13'sd-2937}, {11'sd-963, 12'sd1857, 12'sd1278}, {11'sd-947, 12'sd-1910, 12'sd-1714}},
{{13'sd-2574, 12'sd1886, 11'sd-536}, {12'sd1866, 12'sd1941, 13'sd-2062}, {11'sd-596, 12'sd-1040, 13'sd-2211}},
{{12'sd1373, 13'sd-2421, 10'sd280}, {12'sd-1431, 11'sd907, 12'sd1043}, {12'sd1844, 9'sd-200, 12'sd1420}},
{{13'sd2488, 13'sd-2623, 13'sd-2762}, {13'sd3342, 13'sd2364, 6'sd30}, {12'sd1024, 10'sd508, 12'sd1781}},
{{11'sd643, 12'sd-1742, 11'sd620}, {13'sd2419, 10'sd468, 8'sd-125}, {12'sd1876, 13'sd-2275, 13'sd-2152}},
{{13'sd2415, 12'sd-1917, 13'sd-2967}, {11'sd599, 12'sd-1972, 12'sd-1094}, {7'sd32, 13'sd-2947, 12'sd1176}},
{{13'sd-2527, 12'sd-1281, 12'sd-1027}, {5'sd9, 12'sd2037, 14'sd4677}, {14'sd7993, 14'sd4571, 14'sd4314}},
{{13'sd2331, 13'sd2499, 13'sd2217}, {13'sd-2536, 12'sd1298, 12'sd-1563}, {13'sd-2600, 12'sd-2004, 13'sd-2848}},
{{13'sd-3429, 13'sd-2150, 13'sd2425}, {11'sd-931, 13'sd-2777, 10'sd322}, {11'sd-803, 13'sd-2418, 12'sd1090}},
{{10'sd-481, 11'sd809, 12'sd1148}, {6'sd23, 13'sd2502, 12'sd-1447}, {11'sd-1016, 11'sd-560, 10'sd-312}},
{{12'sd1038, 12'sd-1946, 11'sd635}, {11'sd524, 7'sd-63, 10'sd-281}, {10'sd-475, 11'sd791, 12'sd-1817}},
{{7'sd36, 11'sd785, 12'sd1605}, {12'sd-1310, 7'sd35, 13'sd2962}, {9'sd229, 11'sd641, 12'sd1044}},
{{12'sd1105, 11'sd583, 12'sd-1556}, {10'sd-424, 13'sd-2527, 10'sd-318}, {13'sd-2215, 13'sd-2414, 12'sd-1710}},
{{12'sd-1316, 11'sd-951, 4'sd4}, {12'sd1324, 12'sd-1098, 12'sd1551}, {13'sd-2553, 12'sd-1949, 12'sd1879}},
{{12'sd-1264, 12'sd-1458, 12'sd1130}, {11'sd-575, 12'sd-1856, 6'sd27}, {12'sd1444, 12'sd1790, 11'sd658}},
{{11'sd570, 12'sd1816, 13'sd3333}, {13'sd2468, 11'sd-835, 10'sd-455}, {10'sd-478, 9'sd-226, 13'sd-2960}},
{{10'sd-344, 14'sd-4194, 12'sd-1881}, {12'sd1363, 12'sd1859, 7'sd-51}, {11'sd-938, 11'sd-619, 14'sd4866}},
{{12'sd-1609, 9'sd171, 13'sd-2331}, {12'sd-1865, 13'sd-2350, 8'sd108}, {6'sd17, 12'sd1663, 12'sd1991}},
{{13'sd-2549, 12'sd-1504, 13'sd-2858}, {9'sd-162, 9'sd206, 12'sd1593}, {9'sd235, 12'sd-1860, 13'sd-2352}},
{{13'sd-3177, 13'sd-2747, 6'sd-25}, {1'sd0, 11'sd-714, 13'sd-2261}, {12'sd1887, 12'sd-1539, 11'sd969}},
{{8'sd-70, 11'sd905, 12'sd1396}, {13'sd-3477, 8'sd-108, 10'sd354}, {11'sd880, 13'sd3542, 14'sd4998}},
{{12'sd-1362, 12'sd-1805, 2'sd1}, {11'sd-565, 10'sd390, 13'sd-2128}, {11'sd-921, 13'sd-2566, 13'sd-2586}},
{{11'sd636, 13'sd2460, 9'sd-147}, {13'sd2480, 12'sd1734, 11'sd572}, {12'sd1352, 11'sd-964, 11'sd840}},
{{11'sd913, 11'sd654, 12'sd-1792}, {10'sd472, 7'sd63, 13'sd2771}, {12'sd-1770, 8'sd-82, 12'sd1318}},
{{5'sd8, 8'sd-123, 13'sd2510}, {12'sd-1215, 11'sd-1004, 13'sd-2223}, {7'sd35, 10'sd-432, 14'sd-5875}},
{{12'sd1576, 10'sd-353, 13'sd2895}, {12'sd-1709, 9'sd249, 11'sd-834}, {13'sd2511, 9'sd-132, 13'sd-3103}},
{{14'sd-4388, 12'sd-1331, 13'sd-3684}, {14'sd-5968, 12'sd-1154, 13'sd-3796}, {11'sd-943, 7'sd-50, 5'sd-14}},
{{12'sd1692, 13'sd2514, 12'sd-1584}, {11'sd521, 13'sd2142, 12'sd1899}, {12'sd-1566, 11'sd-723, 12'sd-1785}},
{{12'sd-1670, 12'sd-1941, 12'sd-1781}, {11'sd1000, 10'sd381, 12'sd1562}, {11'sd1008, 12'sd-1937, 13'sd-2466}},
{{12'sd2013, 12'sd-1576, 11'sd-906}, {11'sd1013, 11'sd687, 13'sd-2377}, {5'sd11, 12'sd-1708, 12'sd-1602}},
{{13'sd-3841, 12'sd-1364, 11'sd-537}, {12'sd-1193, 14'sd4418, 11'sd815}, {13'sd2820, 12'sd1508, 13'sd3498}},
{{10'sd353, 13'sd-2681, 12'sd1400}, {12'sd-1110, 11'sd-852, 12'sd-1560}, {12'sd1576, 13'sd2245, 13'sd2204}},
{{12'sd-2037, 12'sd-1133, 12'sd-1542}, {11'sd-559, 12'sd1834, 13'sd-2072}, {9'sd198, 13'sd3388, 8'sd73}},
{{12'sd1121, 12'sd1065, 11'sd996}, {11'sd-584, 12'sd-1144, 12'sd1116}, {12'sd-1121, 10'sd-309, 12'sd-1885}},
{{10'sd336, 13'sd-3041, 13'sd-2799}, {11'sd794, 11'sd-826, 13'sd2503}, {13'sd2435, 12'sd1075, 11'sd975}},
{{13'sd-2331, 12'sd1107, 11'sd-767}, {13'sd3067, 10'sd-457, 12'sd-1566}, {13'sd2317, 13'sd3665, 13'sd2449}},
{{11'sd-518, 11'sd-738, 12'sd1538}, {9'sd-187, 12'sd-1371, 12'sd1790}, {10'sd279, 11'sd583, 13'sd2314}},
{{12'sd1664, 11'sd625, 12'sd-1780}, {11'sd-948, 11'sd-708, 13'sd-2471}, {12'sd-1244, 13'sd2947, 12'sd1834}},
{{13'sd-2514, 12'sd1658, 12'sd-1796}, {13'sd-2084, 11'sd597, 10'sd-454}, {9'sd-204, 9'sd-174, 9'sd-198}},
{{12'sd1492, 12'sd1556, 11'sd907}, {7'sd-41, 11'sd963, 11'sd-995}, {10'sd363, 11'sd-623, 13'sd3256}}},
{
{{13'sd2904, 11'sd879, 8'sd78}, {13'sd2283, 13'sd2804, 13'sd-2519}, {11'sd565, 11'sd696, 13'sd3062}},
{{11'sd828, 13'sd-2064, 10'sd266}, {12'sd1410, 13'sd-2235, 12'sd-1039}, {9'sd210, 13'sd-3232, 12'sd-1642}},
{{13'sd-3186, 12'sd-1751, 13'sd-3265}, {11'sd601, 11'sd662, 12'sd-1921}, {11'sd607, 13'sd2494, 12'sd1291}},
{{12'sd1307, 12'sd1958, 8'sd-92}, {12'sd-1094, 12'sd-1216, 12'sd1533}, {13'sd2082, 10'sd302, 11'sd600}},
{{10'sd293, 12'sd1364, 12'sd1708}, {11'sd813, 13'sd-2799, 13'sd2486}, {13'sd-2505, 6'sd18, 11'sd1005}},
{{7'sd54, 12'sd-1624, 12'sd1270}, {13'sd-2099, 11'sd-571, 7'sd45}, {11'sd803, 11'sd-584, 10'sd-374}},
{{11'sd699, 12'sd-1353, 7'sd-35}, {10'sd306, 11'sd-649, 10'sd281}, {13'sd-3091, 11'sd913, 11'sd614}},
{{11'sd686, 11'sd1017, 13'sd2817}, {12'sd1835, 13'sd-2596, 11'sd-520}, {11'sd-667, 9'sd244, 9'sd-136}},
{{13'sd-2968, 12'sd1674, 12'sd1041}, {12'sd-1229, 12'sd-1471, 13'sd2305}, {9'sd-229, 9'sd193, 12'sd1417}},
{{12'sd1756, 13'sd2229, 13'sd2580}, {12'sd1786, 13'sd2296, 11'sd-637}, {11'sd1005, 12'sd1362, 11'sd-839}},
{{13'sd-2582, 9'sd213, 12'sd-1854}, {12'sd-1721, 12'sd1681, 13'sd2062}, {13'sd2207, 11'sd-882, 11'sd784}},
{{11'sd1004, 13'sd2401, 12'sd1837}, {13'sd2383, 13'sd2396, 12'sd1388}, {11'sd-815, 12'sd-1536, 12'sd1323}},
{{11'sd-552, 7'sd-43, 13'sd2804}, {12'sd1398, 10'sd279, 13'sd2297}, {10'sd-507, 13'sd2899, 12'sd1100}},
{{9'sd209, 12'sd-1936, 13'sd2414}, {12'sd-1397, 10'sd-302, 12'sd-1194}, {13'sd-2603, 10'sd-261, 8'sd-73}},
{{13'sd-3178, 10'sd270, 12'sd1894}, {9'sd-215, 10'sd263, 11'sd-1016}, {13'sd2467, 13'sd-2198, 11'sd-956}},
{{12'sd1640, 11'sd557, 11'sd764}, {9'sd-166, 11'sd-857, 12'sd1369}, {11'sd-588, 13'sd2065, 5'sd15}},
{{11'sd-889, 13'sd-2692, 12'sd-1280}, {12'sd-1734, 13'sd-2131, 10'sd316}, {13'sd-2419, 12'sd1996, 13'sd2116}},
{{9'sd250, 12'sd1177, 11'sd998}, {12'sd1167, 13'sd2875, 13'sd2412}, {10'sd479, 13'sd3819, 13'sd3782}},
{{13'sd-2856, 11'sd-578, 13'sd2857}, {12'sd1088, 9'sd209, 11'sd648}, {12'sd1944, 12'sd-1713, 12'sd1272}},
{{13'sd-2392, 12'sd1117, 11'sd790}, {12'sd1236, 10'sd-487, 13'sd2474}, {6'sd-27, 12'sd-1430, 13'sd-2055}},
{{13'sd2248, 13'sd2968, 13'sd-2870}, {12'sd-2013, 12'sd-1963, 10'sd357}, {11'sd-1010, 9'sd-247, 11'sd959}},
{{8'sd77, 12'sd-1082, 12'sd1524}, {6'sd-31, 11'sd-919, 12'sd-1432}, {12'sd1747, 11'sd964, 12'sd-1490}},
{{12'sd-1462, 13'sd-3047, 11'sd837}, {13'sd2193, 13'sd-2338, 12'sd1468}, {11'sd810, 9'sd212, 13'sd2663}},
{{11'sd-617, 13'sd2210, 6'sd-19}, {10'sd316, 10'sd-375, 13'sd2839}, {10'sd-477, 13'sd-3134, 13'sd2378}},
{{12'sd-1399, 11'sd-820, 13'sd-3011}, {10'sd487, 11'sd-539, 13'sd-2088}, {13'sd2095, 13'sd2434, 13'sd2201}},
{{12'sd1759, 13'sd-2270, 12'sd1441}, {10'sd322, 13'sd2325, 12'sd-1148}, {12'sd1167, 13'sd2143, 12'sd-1266}},
{{12'sd1301, 9'sd137, 9'sd-138}, {12'sd1877, 12'sd-1253, 10'sd-291}, {13'sd2333, 9'sd-245, 11'sd914}},
{{12'sd-1090, 10'sd311, 11'sd904}, {12'sd1458, 12'sd1332, 11'sd916}, {13'sd-2165, 11'sd-990, 12'sd1233}},
{{12'sd-1840, 10'sd321, 8'sd71}, {11'sd756, 13'sd2237, 11'sd987}, {13'sd2866, 10'sd-361, 11'sd988}},
{{12'sd1481, 13'sd-2122, 9'sd195}, {13'sd-2382, 11'sd-815, 13'sd-2475}, {8'sd-111, 13'sd-2811, 11'sd-897}},
{{11'sd-648, 12'sd1322, 13'sd2190}, {12'sd-1711, 11'sd-637, 12'sd1830}, {11'sd-785, 13'sd-2576, 11'sd1009}},
{{12'sd1686, 10'sd403, 11'sd-902}, {13'sd2223, 12'sd-1610, 10'sd306}, {11'sd-514, 13'sd2818, 11'sd721}},
{{10'sd398, 12'sd-1939, 11'sd-918}, {13'sd3677, 11'sd-754, 13'sd2620}, {13'sd3053, 13'sd2526, 12'sd1929}},
{{14'sd-4615, 12'sd1525, 11'sd-905}, {11'sd858, 13'sd2295, 11'sd611}, {13'sd-2294, 12'sd-1582, 13'sd-2156}},
{{12'sd-1727, 13'sd-2252, 11'sd985}, {12'sd-1642, 12'sd1908, 12'sd1715}, {12'sd-1173, 12'sd-1229, 13'sd-2605}},
{{13'sd-2505, 13'sd2440, 11'sd727}, {12'sd1705, 9'sd158, 12'sd-1776}, {12'sd-1522, 12'sd-1278, 12'sd-1738}},
{{12'sd1669, 12'sd-1636, 12'sd-1371}, {11'sd769, 11'sd692, 12'sd1416}, {12'sd-1230, 12'sd1137, 12'sd-1730}},
{{12'sd-1457, 11'sd-656, 12'sd-1117}, {11'sd-691, 12'sd-1029, 12'sd1952}, {12'sd-1579, 13'sd-2581, 7'sd-55}},
{{12'sd-1123, 11'sd820, 12'sd1481}, {9'sd151, 12'sd1548, 11'sd798}, {10'sd-348, 12'sd1746, 12'sd-1644}},
{{11'sd687, 11'sd-817, 12'sd1315}, {12'sd-1480, 13'sd-2258, 11'sd-792}, {9'sd-183, 12'sd-1425, 11'sd-826}},
{{13'sd3018, 10'sd-397, 13'sd3262}, {11'sd866, 13'sd2987, 13'sd3393}, {14'sd4310, 11'sd973, 10'sd497}},
{{9'sd-165, 11'sd-860, 11'sd-645}, {13'sd2873, 12'sd-1375, 12'sd-1662}, {13'sd2813, 13'sd3800, 12'sd-1574}},
{{11'sd-1016, 13'sd-3296, 12'sd-1396}, {9'sd166, 12'sd1441, 12'sd-1344}, {12'sd-1676, 13'sd3007, 13'sd2082}},
{{11'sd-523, 10'sd329, 13'sd2575}, {12'sd-1049, 8'sd-90, 13'sd2599}, {13'sd2740, 12'sd1173, 9'sd-203}},
{{13'sd-3929, 12'sd1613, 9'sd204}, {11'sd-943, 13'sd-2423, 12'sd1665}, {11'sd-960, 13'sd2231, 12'sd1638}},
{{13'sd-2283, 10'sd459, 10'sd-367}, {12'sd-1742, 11'sd-527, 12'sd1884}, {11'sd-826, 11'sd575, 11'sd1007}},
{{12'sd-1966, 11'sd764, 12'sd1673}, {11'sd746, 13'sd2841, 13'sd2302}, {12'sd-1836, 11'sd-860, 13'sd2745}},
{{12'sd-1344, 13'sd-2372, 11'sd-591}, {12'sd-1122, 7'sd49, 13'sd2247}, {6'sd-21, 11'sd659, 12'sd1423}},
{{13'sd2181, 13'sd3544, 11'sd-689}, {11'sd832, 10'sd-415, 12'sd-1408}, {13'sd-2636, 13'sd3145, 13'sd2160}},
{{13'sd3168, 12'sd1294, 14'sd5274}, {13'sd2695, 9'sd251, 13'sd2436}, {11'sd-642, 11'sd934, 13'sd4035}},
{{6'sd31, 8'sd110, 12'sd-1126}, {12'sd1257, 11'sd-888, 14'sd-4274}, {12'sd1839, 11'sd-679, 11'sd-686}},
{{12'sd-1053, 13'sd2933, 13'sd2448}, {12'sd1643, 11'sd861, 9'sd178}, {12'sd1424, 9'sd-230, 13'sd-2278}},
{{13'sd-2571, 13'sd-2422, 12'sd-1586}, {12'sd1913, 12'sd1720, 10'sd391}, {13'sd-2098, 12'sd1687, 12'sd1689}},
{{12'sd-1566, 12'sd1639, 11'sd697}, {12'sd-1156, 12'sd-1382, 12'sd1497}, {11'sd581, 13'sd-2636, 13'sd-3291}},
{{12'sd-1510, 11'sd920, 9'sd-182}, {12'sd1125, 12'sd1687, 13'sd-2068}, {14'sd5543, 12'sd1160, 13'sd2358}},
{{12'sd-1629, 13'sd-2303, 9'sd206}, {13'sd-2674, 11'sd-609, 11'sd906}, {11'sd-975, 12'sd1371, 13'sd2197}},
{{12'sd-1274, 12'sd1260, 12'sd-1305}, {11'sd-702, 12'sd-1791, 11'sd-865}, {13'sd2123, 12'sd-1213, 10'sd-374}},
{{9'sd255, 9'sd-182, 11'sd632}, {9'sd131, 13'sd-2400, 11'sd-561}, {11'sd-650, 13'sd-3251, 5'sd8}},
{{13'sd-2085, 6'sd16, 12'sd-1891}, {11'sd887, 9'sd251, 11'sd-909}, {14'sd-4437, 10'sd407, 13'sd-3172}},
{{5'sd-11, 10'sd-387, 14'sd-4390}, {11'sd975, 10'sd425, 13'sd-2571}, {10'sd419, 13'sd2402, 12'sd-1919}},
{{13'sd-2563, 10'sd292, 8'sd93}, {12'sd1489, 12'sd1025, 13'sd-2226}, {11'sd-557, 12'sd1705, 13'sd-2165}},
{{13'sd3845, 13'sd2544, 12'sd1625}, {12'sd1568, 12'sd1729, 13'sd2584}, {11'sd806, 12'sd1673, 13'sd-2793}},
{{9'sd147, 6'sd-31, 13'sd-2091}, {13'sd2482, 13'sd-2313, 13'sd-3968}, {11'sd1006, 12'sd-1873, 10'sd460}},
{{12'sd1394, 12'sd-1453, 11'sd583}, {12'sd1661, 11'sd-843, 13'sd3300}, {10'sd-454, 10'sd-474, 13'sd2651}}},
{
{{9'sd-233, 12'sd-1551, 11'sd908}, {13'sd2459, 12'sd1138, 12'sd-1162}, {6'sd24, 12'sd-1164, 12'sd-1137}},
{{11'sd-983, 12'sd1454, 12'sd1931}, {13'sd-2327, 11'sd800, 13'sd-2656}, {10'sd429, 13'sd-2143, 12'sd1977}},
{{13'sd2818, 13'sd3326, 13'sd4013}, {9'sd-151, 13'sd-2136, 10'sd443}, {12'sd-1361, 14'sd-4457, 7'sd-59}},
{{11'sd584, 12'sd-1719, 12'sd-1959}, {11'sd597, 13'sd-3506, 13'sd-2716}, {11'sd680, 12'sd-1228, 8'sd-90}},
{{6'sd-18, 10'sd-263, 12'sd1670}, {12'sd1257, 10'sd-509, 10'sd-454}, {12'sd-1815, 12'sd1108, 11'sd682}},
{{8'sd83, 11'sd907, 12'sd1714}, {13'sd-2306, 12'sd-1083, 13'sd-2505}, {12'sd-1184, 12'sd1566, 12'sd1234}},
{{10'sd-282, 13'sd-2301, 11'sd525}, {11'sd-880, 11'sd839, 13'sd-2833}, {9'sd-234, 11'sd615, 11'sd868}},
{{11'sd-727, 12'sd1370, 11'sd-958}, {12'sd-1136, 9'sd-165, 13'sd-2081}, {6'sd17, 13'sd-2499, 12'sd-1650}},
{{12'sd-1120, 10'sd297, 12'sd-1925}, {12'sd-1100, 12'sd-1669, 10'sd-494}, {10'sd496, 13'sd-3237, 11'sd-626}},
{{12'sd-2037, 11'sd-630, 12'sd-1386}, {12'sd-1904, 11'sd769, 11'sd595}, {11'sd-982, 12'sd1411, 12'sd-1735}},
{{8'sd127, 13'sd-3017, 11'sd-598}, {13'sd-2694, 13'sd-2792, 12'sd-1278}, {12'sd-1950, 11'sd-580, 11'sd588}},
{{11'sd-1017, 11'sd949, 12'sd1381}, {11'sd-1001, 12'sd-1749, 12'sd1563}, {12'sd1621, 12'sd-1894, 10'sd476}},
{{12'sd-1794, 13'sd-3501, 13'sd-2846}, {11'sd902, 11'sd-558, 13'sd-2947}, {12'sd1033, 13'sd-2412, 13'sd-3075}},
{{11'sd748, 12'sd-1412, 13'sd2272}, {12'sd-1569, 12'sd1116, 12'sd2012}, {13'sd2754, 9'sd246, 13'sd-2646}},
{{12'sd-1547, 12'sd1538, 12'sd1031}, {12'sd1372, 13'sd2373, 12'sd-1403}, {13'sd-2910, 12'sd1046, 9'sd163}},
{{11'sd-1021, 12'sd2008, 12'sd1591}, {12'sd2047, 12'sd1274, 12'sd-1080}, {12'sd1637, 12'sd1326, 11'sd-583}},
{{12'sd1899, 12'sd1337, 7'sd-42}, {12'sd1578, 11'sd624, 11'sd-702}, {11'sd-513, 13'sd2832, 11'sd680}},
{{13'sd2445, 8'sd77, 11'sd-894}, {10'sd-304, 11'sd650, 9'sd144}, {13'sd-2547, 12'sd1229, 10'sd303}},
{{13'sd2464, 12'sd-1590, 11'sd577}, {13'sd2204, 13'sd-2230, 10'sd302}, {12'sd-1796, 11'sd-555, 12'sd-2011}},
{{12'sd-1111, 12'sd-1088, 13'sd-2052}, {11'sd694, 9'sd-140, 13'sd-2645}, {13'sd2409, 13'sd-2554, 12'sd-1571}},
{{11'sd521, 7'sd50, 12'sd2004}, {13'sd-2835, 12'sd1260, 11'sd-727}, {12'sd1535, 13'sd2175, 12'sd1281}},
{{12'sd1578, 11'sd798, 11'sd-947}, {13'sd2110, 13'sd-3394, 9'sd-130}, {12'sd-1556, 12'sd-1498, 12'sd-1492}},
{{13'sd2138, 12'sd-1442, 12'sd1076}, {12'sd1312, 13'sd2171, 10'sd-356}, {12'sd-1336, 12'sd1851, 12'sd1326}},
{{10'sd-431, 12'sd-1546, 13'sd2429}, {10'sd-304, 13'sd2635, 11'sd520}, {13'sd2871, 12'sd-1146, 12'sd1608}},
{{11'sd-670, 13'sd-2140, 13'sd2083}, {12'sd-1754, 12'sd1425, 12'sd1914}, {12'sd1933, 11'sd-978, 12'sd1280}},
{{11'sd605, 11'sd558, 9'sd-147}, {10'sd-333, 10'sd-278, 10'sd-456}, {12'sd1761, 11'sd-661, 13'sd-2114}},
{{11'sd-862, 12'sd-1801, 12'sd1343}, {12'sd1503, 12'sd-1927, 11'sd864}, {10'sd273, 12'sd1957, 11'sd937}},
{{11'sd-787, 13'sd-2312, 13'sd-2749}, {12'sd1231, 9'sd-133, 13'sd-2327}, {11'sd524, 9'sd-172, 12'sd1512}},
{{13'sd-2170, 12'sd-1807, 13'sd2881}, {9'sd239, 11'sd-911, 13'sd2910}, {13'sd-2849, 13'sd-3420, 12'sd-1126}},
{{13'sd-3368, 12'sd1437, 13'sd-2858}, {10'sd-477, 12'sd-1258, 11'sd749}, {12'sd-1058, 13'sd-2169, 5'sd-12}},
{{12'sd-1322, 13'sd3147, 12'sd1730}, {12'sd1656, 13'sd3336, 12'sd-1100}, {11'sd-635, 12'sd1571, 12'sd1152}},
{{12'sd1540, 13'sd2432, 11'sd802}, {9'sd-164, 12'sd1234, 12'sd-1376}, {12'sd-1092, 12'sd-1365, 12'sd1200}},
{{13'sd-3502, 13'sd-2658, 11'sd-565}, {10'sd372, 12'sd1610, 13'sd3120}, {12'sd-1477, 12'sd1877, 13'sd3385}},
{{11'sd-844, 11'sd709, 11'sd962}, {9'sd141, 13'sd2565, 12'sd1104}, {13'sd-2598, 13'sd-2721, 11'sd534}},
{{12'sd-1926, 13'sd-2672, 11'sd545}, {11'sd-996, 12'sd-1573, 12'sd1581}, {13'sd-3015, 13'sd-3162, 11'sd914}},
{{11'sd811, 11'sd-639, 10'sd304}, {12'sd-1518, 9'sd143, 12'sd1094}, {13'sd-2828, 12'sd1298, 12'sd-1736}},
{{13'sd-2426, 13'sd-2293, 10'sd343}, {11'sd879, 12'sd1451, 11'sd954}, {11'sd891, 12'sd1432, 13'sd-2472}},
{{12'sd-1465, 12'sd-1345, 13'sd-2165}, {11'sd628, 13'sd2641, 10'sd302}, {13'sd2236, 13'sd-2179, 12'sd-1525}},
{{12'sd1682, 12'sd-1217, 13'sd-2462}, {13'sd2455, 11'sd522, 10'sd415}, {12'sd1271, 13'sd2508, 12'sd-1115}},
{{12'sd1298, 12'sd1417, 13'sd-2865}, {9'sd-183, 9'sd249, 11'sd-859}, {8'sd-66, 12'sd1821, 12'sd1695}},
{{13'sd2810, 12'sd-1691, 13'sd-4006}, {12'sd1763, 12'sd-1498, 11'sd785}, {10'sd-372, 12'sd-1262, 12'sd1099}},
{{12'sd1594, 12'sd1111, 12'sd1334}, {11'sd-542, 13'sd-3481, 13'sd2435}, {13'sd-2979, 12'sd-1624, 13'sd-3797}},
{{13'sd-2057, 12'sd1770, 13'sd2770}, {9'sd225, 12'sd-1286, 10'sd434}, {13'sd-2557, 9'sd-164, 12'sd1535}},
{{11'sd-941, 13'sd2266, 12'sd-1502}, {12'sd1692, 11'sd-737, 10'sd280}, {12'sd1075, 12'sd-1712, 4'sd-5}},
{{13'sd3100, 9'sd-225, 12'sd1431}, {11'sd-953, 13'sd-2671, 12'sd-1602}, {9'sd-152, 9'sd-218, 13'sd-3531}},
{{13'sd-2655, 12'sd-1483, 11'sd941}, {10'sd281, 8'sd107, 13'sd-2812}, {7'sd-35, 13'sd2568, 12'sd1726}},
{{11'sd605, 12'sd1793, 13'sd2287}, {13'sd-2863, 10'sd353, 13'sd-2519}, {12'sd-1793, 10'sd-265, 12'sd1322}},
{{11'sd945, 11'sd-631, 11'sd-930}, {12'sd-1235, 13'sd2125, 12'sd-1384}, {12'sd-1684, 12'sd-1452, 12'sd-1851}},
{{10'sd-405, 12'sd-1168, 12'sd1677}, {13'sd2646, 13'sd3103, 12'sd1636}, {13'sd-2120, 13'sd2703, 12'sd2004}},
{{13'sd-2377, 12'sd-1587, 13'sd-3073}, {13'sd2686, 12'sd1776, 12'sd-1703}, {12'sd1981, 13'sd2130, 10'sd389}},
{{13'sd2192, 11'sd612, 13'sd3605}, {11'sd706, 13'sd2945, 11'sd781}, {11'sd599, 10'sd385, 12'sd-1341}},
{{11'sd723, 10'sd-471, 13'sd-2874}, {13'sd2351, 13'sd-2939, 11'sd-792}, {12'sd-1444, 13'sd-3353, 12'sd-1242}},
{{12'sd-1883, 12'sd1370, 12'sd1045}, {12'sd1036, 10'sd-260, 11'sd762}, {12'sd-1653, 7'sd57, 11'sd-808}},
{{8'sd-96, 11'sd694, 11'sd642}, {13'sd-2542, 12'sd1377, 12'sd1700}, {11'sd784, 13'sd2060, 13'sd3128}},
{{11'sd-979, 13'sd3381, 13'sd3748}, {13'sd-3548, 13'sd-2813, 12'sd1264}, {14'sd-4828, 14'sd-4293, 12'sd1926}},
{{11'sd-909, 11'sd-611, 13'sd2420}, {10'sd267, 13'sd-2188, 12'sd-1843}, {12'sd-1971, 12'sd-1127, 10'sd-336}},
{{12'sd-1522, 11'sd657, 12'sd-1553}, {13'sd-2670, 11'sd-552, 11'sd602}, {13'sd-3186, 13'sd-3411, 12'sd-2032}},
{{12'sd-1770, 13'sd2390, 12'sd-1307}, {12'sd1547, 12'sd1473, 11'sd-670}, {11'sd-601, 13'sd2391, 13'sd-2939}},
{{13'sd-3095, 7'sd60, 13'sd2637}, {12'sd1960, 12'sd1795, 12'sd1237}, {12'sd-1441, 11'sd693, 10'sd-269}},
{{10'sd-498, 13'sd-2169, 12'sd1180}, {12'sd-1701, 13'sd-2204, 13'sd-3045}, {10'sd475, 12'sd-2004, 13'sd-2537}},
{{12'sd1760, 12'sd1705, 11'sd-827}, {11'sd705, 11'sd-936, 9'sd-176}, {13'sd2691, 10'sd-404, 11'sd999}},
{{12'sd1171, 10'sd383, 11'sd-819}, {8'sd-87, 11'sd724, 11'sd-552}, {12'sd1466, 11'sd799, 8'sd-89}},
{{12'sd1314, 7'sd-35, 11'sd853}, {9'sd-218, 13'sd2319, 12'sd1554}, {10'sd-261, 13'sd-2201, 13'sd2247}},
{{13'sd3455, 13'sd3430, 11'sd923}, {12'sd-1646, 12'sd1421, 10'sd305}, {12'sd-1240, 13'sd2179, 13'sd-2593}}},
{
{{11'sd-874, 11'sd990, 11'sd-1012}, {12'sd-1449, 13'sd2095, 13'sd-2117}, {9'sd-255, 11'sd808, 12'sd-1253}},
{{13'sd2438, 13'sd-2324, 13'sd2455}, {12'sd2037, 10'sd464, 13'sd2952}, {7'sd46, 12'sd-1396, 12'sd1558}},
{{14'sd-4681, 8'sd92, 9'sd156}, {9'sd-172, 12'sd1580, 13'sd2100}, {11'sd776, 13'sd-3700, 12'sd-1743}},
{{11'sd890, 10'sd-479, 10'sd-334}, {10'sd322, 13'sd-2355, 11'sd-788}, {10'sd498, 12'sd-1813, 12'sd-2013}},
{{10'sd458, 11'sd789, 11'sd-782}, {12'sd2024, 12'sd-1482, 13'sd-2098}, {13'sd-2277, 13'sd2554, 10'sd357}},
{{11'sd725, 13'sd-2491, 12'sd1691}, {13'sd2203, 11'sd609, 12'sd-1452}, {13'sd2845, 10'sd-277, 12'sd-1156}},
{{12'sd-1054, 12'sd1318, 12'sd1479}, {12'sd-1542, 11'sd731, 13'sd3111}, {11'sd-1000, 10'sd-323, 12'sd1730}},
{{12'sd1645, 10'sd331, 12'sd1369}, {13'sd2052, 11'sd993, 12'sd-1780}, {12'sd-1815, 13'sd-2085, 11'sd860}},
{{12'sd-1924, 13'sd-2676, 13'sd-3537}, {11'sd-555, 13'sd-2318, 9'sd212}, {10'sd310, 13'sd-2403, 12'sd-1771}},
{{13'sd2450, 11'sd514, 11'sd-814}, {10'sd-431, 12'sd-1075, 9'sd171}, {9'sd-175, 4'sd4, 13'sd2097}},
{{13'sd2359, 12'sd-1828, 13'sd2349}, {10'sd-364, 12'sd-1038, 13'sd3215}, {11'sd-517, 11'sd631, 13'sd2183}},
{{11'sd941, 12'sd-1955, 9'sd160}, {13'sd3011, 11'sd571, 13'sd2480}, {12'sd2000, 7'sd54, 12'sd-1789}},
{{11'sd694, 14'sd-4097, 14'sd-4760}, {13'sd2535, 11'sd530, 12'sd2037}, {11'sd654, 12'sd1088, 11'sd553}},
{{9'sd-187, 6'sd26, 13'sd2455}, {10'sd-389, 12'sd-2008, 12'sd1390}, {11'sd-773, 12'sd-1585, 10'sd-405}},
{{11'sd755, 12'sd1292, 13'sd-2895}, {10'sd334, 13'sd-2189, 10'sd-500}, {12'sd1159, 11'sd674, 8'sd-98}},
{{11'sd-1023, 13'sd2406, 13'sd2088}, {13'sd-2375, 11'sd-868, 12'sd-1348}, {12'sd1371, 13'sd2500, 13'sd3047}},
{{12'sd1092, 12'sd-1211, 10'sd284}, {12'sd-1158, 11'sd-767, 13'sd-2310}, {12'sd-2011, 11'sd720, 12'sd1590}},
{{11'sd642, 13'sd2974, 12'sd1969}, {11'sd-771, 11'sd1002, 12'sd-1569}, {14'sd-5447, 13'sd-2350, 13'sd-3100}},
{{13'sd-2152, 13'sd2097, 13'sd2199}, {13'sd-2494, 12'sd-1086, 12'sd1253}, {12'sd-1840, 12'sd1105, 10'sd378}},
{{12'sd1531, 9'sd222, 13'sd2989}, {11'sd941, 12'sd1925, 11'sd-1022}, {12'sd-1697, 12'sd1464, 13'sd2571}},
{{12'sd1422, 12'sd-1712, 9'sd-148}, {13'sd2973, 11'sd-960, 10'sd416}, {10'sd-318, 11'sd1023, 12'sd1602}},
{{12'sd-1779, 10'sd457, 13'sd-3197}, {12'sd1773, 12'sd-1639, 13'sd2244}, {13'sd-2298, 12'sd-1237, 12'sd-1702}},
{{12'sd1187, 11'sd-581, 11'sd835}, {10'sd-382, 11'sd-887, 10'sd-404}, {12'sd1196, 11'sd-800, 12'sd-1187}},
{{13'sd-2152, 11'sd531, 13'sd3022}, {11'sd941, 6'sd18, 13'sd2113}, {11'sd-668, 11'sd838, 12'sd1516}},
{{13'sd-2067, 12'sd-1838, 13'sd-2186}, {13'sd2838, 12'sd-1689, 13'sd-2279}, {13'sd2868, 11'sd-929, 10'sd497}},
{{12'sd1565, 13'sd2092, 12'sd1512}, {12'sd1668, 5'sd-11, 12'sd-1761}, {10'sd-427, 13'sd-2471, 12'sd1353}},
{{12'sd-1291, 12'sd1205, 13'sd-2243}, {8'sd-83, 12'sd-1954, 12'sd1394}, {11'sd803, 12'sd1534, 12'sd-1051}},
{{13'sd2207, 12'sd1376, 13'sd-2160}, {12'sd1269, 13'sd2442, 11'sd-667}, {13'sd3334, 9'sd155, 13'sd2514}},
{{12'sd1725, 13'sd-2858, 12'sd-1540}, {12'sd2033, 6'sd24, 13'sd-2183}, {12'sd1210, 12'sd1411, 10'sd364}},
{{11'sd717, 12'sd-1323, 12'sd-1736}, {7'sd39, 5'sd-15, 13'sd-2587}, {11'sd-793, 12'sd-1265, 11'sd1005}},
{{13'sd3637, 11'sd647, 13'sd2412}, {13'sd2084, 13'sd2486, 12'sd1172}, {12'sd1404, 13'sd2487, 13'sd3067}},
{{9'sd-197, 13'sd-2647, 12'sd1911}, {12'sd1841, 12'sd1729, 10'sd443}, {12'sd1339, 11'sd-735, 11'sd678}},
{{11'sd-851, 11'sd-971, 12'sd-1834}, {13'sd2196, 12'sd1514, 13'sd2595}, {10'sd358, 13'sd3695, 13'sd2219}},
{{11'sd798, 10'sd403, 12'sd1035}, {13'sd2742, 13'sd2601, 10'sd365}, {12'sd-1934, 11'sd766, 10'sd-258}},
{{12'sd-1732, 11'sd673, 13'sd-2645}, {13'sd2722, 13'sd2563, 12'sd1269}, {11'sd616, 12'sd1071, 11'sd-989}},
{{13'sd-2056, 13'sd2292, 1'sd0}, {11'sd845, 11'sd812, 12'sd1610}, {12'sd1210, 11'sd655, 12'sd-1241}},
{{13'sd-2419, 9'sd141, 12'sd-1060}, {12'sd1057, 9'sd-224, 13'sd2760}, {9'sd-183, 12'sd1841, 13'sd2996}},
{{12'sd-1704, 10'sd423, 12'sd-1091}, {13'sd2509, 13'sd2069, 10'sd461}, {12'sd1383, 12'sd-1646, 11'sd746}},
{{13'sd3869, 12'sd1321, 13'sd2513}, {13'sd3533, 12'sd-1493, 6'sd-24}, {8'sd-96, 11'sd-575, 12'sd1480}},
{{12'sd1193, 11'sd-541, 13'sd2857}, {11'sd-995, 12'sd2027, 12'sd1639}, {13'sd2751, 13'sd2141, 13'sd3430}},
{{13'sd-3091, 11'sd-916, 13'sd-2754}, {13'sd-3263, 10'sd368, 7'sd-61}, {12'sd1360, 10'sd435, 13'sd2226}},
{{12'sd-1172, 13'sd-2416, 13'sd-3904}, {11'sd-725, 7'sd-50, 13'sd-2637}, {12'sd1084, 13'sd-2106, 12'sd-2000}},
{{11'sd576, 12'sd-1124, 12'sd2016}, {12'sd1832, 13'sd2507, 13'sd2590}, {11'sd559, 13'sd-2322, 13'sd2435}},
{{13'sd-2280, 13'sd2761, 12'sd1256}, {12'sd-1781, 10'sd456, 12'sd1354}, {13'sd-2728, 11'sd-630, 12'sd1316}},
{{12'sd-1838, 13'sd-2593, 9'sd237}, {12'sd1574, 7'sd-48, 11'sd806}, {12'sd2046, 12'sd1382, 12'sd1384}},
{{12'sd1775, 11'sd577, 9'sd-161}, {12'sd-1440, 12'sd1312, 12'sd-1383}, {12'sd1600, 9'sd156, 12'sd-1053}},
{{13'sd-2115, 11'sd-876, 8'sd78}, {9'sd230, 12'sd1364, 13'sd-2066}, {10'sd-350, 12'sd-1506, 10'sd409}},
{{13'sd-2308, 10'sd345, 12'sd-1593}, {9'sd201, 13'sd-2316, 10'sd314}, {13'sd-2324, 12'sd1385, 8'sd105}},
{{12'sd-1515, 9'sd191, 13'sd2293}, {12'sd-1092, 12'sd-1867, 13'sd2402}, {13'sd-2873, 12'sd1678, 14'sd4202}},
{{13'sd-2767, 12'sd1523, 12'sd1112}, {8'sd-116, 13'sd-2124, 11'sd-638}, {12'sd1438, 13'sd3331, 11'sd557}},
{{12'sd-1389, 13'sd-2540, 9'sd-130}, {12'sd1722, 9'sd-210, 12'sd1377}, {12'sd2046, 8'sd99, 11'sd-673}},
{{12'sd1462, 13'sd-2927, 13'sd-2261}, {13'sd-2111, 13'sd2074, 12'sd-1244}, {13'sd-2171, 12'sd1249, 11'sd-696}},
{{11'sd-975, 9'sd-218, 11'sd694}, {13'sd2891, 12'sd1323, 13'sd2397}, {10'sd-379, 13'sd2958, 12'sd1070}},
{{9'sd145, 13'sd-2085, 13'sd-2343}, {13'sd-2561, 12'sd-1499, 8'sd81}, {3'sd2, 12'sd1892, 10'sd-279}},
{{13'sd2076, 11'sd761, 12'sd-1543}, {13'sd2684, 10'sd-371, 11'sd951}, {8'sd71, 13'sd-2972, 12'sd-1554}},
{{12'sd1283, 12'sd2007, 13'sd-2717}, {12'sd1561, 13'sd2841, 13'sd-2711}, {11'sd-610, 10'sd344, 12'sd-1939}},
{{10'sd-310, 13'sd2065, 13'sd2434}, {12'sd-1540, 11'sd912, 11'sd891}, {11'sd-542, 10'sd-421, 12'sd-1141}},
{{10'sd-509, 12'sd-1641, 12'sd-1964}, {12'sd1836, 13'sd3404, 11'sd652}, {11'sd-525, 12'sd-1387, 12'sd1804}},
{{12'sd1195, 6'sd23, 13'sd3255}, {12'sd1676, 12'sd1877, 11'sd-1007}, {8'sd-66, 12'sd-1613, 12'sd1186}},
{{13'sd2492, 9'sd144, 12'sd-1228}, {12'sd1220, 11'sd-515, 12'sd-1640}, {13'sd-2332, 13'sd-3826, 11'sd-528}},
{{13'sd-2310, 13'sd2555, 9'sd-134}, {11'sd-924, 12'sd2015, 8'sd125}, {12'sd-1107, 11'sd655, 12'sd-1669}},
{{9'sd-211, 13'sd2084, 11'sd-843}, {10'sd329, 13'sd2156, 13'sd2612}, {12'sd-1977, 10'sd-340, 8'sd119}},
{{12'sd-1406, 11'sd-1005, 11'sd532}, {12'sd1904, 13'sd2330, 13'sd-2170}, {13'sd2207, 11'sd808, 13'sd2082}},
{{12'sd1135, 13'sd-2546, 11'sd878}, {11'sd587, 12'sd1585, 10'sd369}, {13'sd-2685, 13'sd-2364, 13'sd-2402}}},
{
{{6'sd18, 11'sd965, 8'sd-85}, {13'sd-3972, 12'sd-1514, 12'sd1260}, {10'sd-352, 12'sd1635, 13'sd-2071}},
{{12'sd-1117, 11'sd734, 12'sd-1804}, {12'sd-1285, 12'sd1200, 12'sd1457}, {10'sd403, 11'sd860, 13'sd2741}},
{{14'sd4583, 13'sd3008, 10'sd371}, {12'sd-1139, 12'sd1770, 12'sd1347}, {12'sd1778, 12'sd1515, 12'sd-1180}},
{{12'sd1111, 13'sd2546, 4'sd-4}, {12'sd-1388, 13'sd-2184, 12'sd-1708}, {13'sd-2929, 12'sd1323, 13'sd-2971}},
{{10'sd288, 12'sd-1470, 12'sd1625}, {13'sd2070, 13'sd2716, 11'sd-649}, {10'sd-435, 13'sd2763, 13'sd-2140}},
{{13'sd-2711, 13'sd2706, 12'sd1082}, {13'sd-3085, 12'sd1392, 12'sd1045}, {12'sd-1756, 8'sd105, 8'sd-99}},
{{13'sd-3746, 13'sd-2578, 9'sd-131}, {12'sd-1058, 12'sd1465, 12'sd-1617}, {12'sd1786, 12'sd-1419, 11'sd968}},
{{12'sd1707, 12'sd-1092, 11'sd754}, {12'sd1153, 9'sd173, 11'sd655}, {11'sd953, 11'sd-984, 12'sd1128}},
{{11'sd986, 12'sd1602, 12'sd1084}, {14'sd4171, 13'sd-2051, 13'sd2901}, {13'sd-2741, 12'sd-1790, 12'sd1303}},
{{13'sd-2839, 13'sd-2202, 9'sd-236}, {10'sd425, 11'sd778, 12'sd-1160}, {13'sd-3221, 12'sd-1233, 12'sd-1555}},
{{13'sd3047, 12'sd-1919, 12'sd-1958}, {12'sd-1034, 11'sd624, 12'sd-1942}, {13'sd2142, 8'sd95, 12'sd1667}},
{{11'sd572, 13'sd3415, 12'sd-1478}, {12'sd1151, 9'sd-226, 12'sd1276}, {13'sd-2346, 13'sd2383, 10'sd508}},
{{9'sd157, 12'sd1874, 12'sd1613}, {6'sd19, 11'sd660, 9'sd-175}, {12'sd-1103, 11'sd-792, 10'sd454}},
{{10'sd457, 12'sd-1223, 13'sd-2330}, {13'sd-3375, 13'sd-2455, 12'sd-1451}, {12'sd-1091, 8'sd-80, 12'sd1223}},
{{12'sd1221, 13'sd2931, 14'sd4664}, {10'sd-374, 12'sd-1864, 13'sd4075}, {12'sd-1179, 12'sd2044, 14'sd4999}},
{{12'sd-1202, 12'sd-1881, 9'sd129}, {11'sd-777, 12'sd1672, 12'sd1581}, {13'sd-3811, 12'sd-1620, 10'sd270}},
{{13'sd-2586, 13'sd-2738, 12'sd-1913}, {13'sd-2425, 12'sd1822, 10'sd413}, {12'sd1276, 12'sd1857, 12'sd1827}},
{{11'sd-1010, 13'sd3036, 9'sd140}, {12'sd1181, 11'sd-871, 12'sd-1447}, {12'sd1449, 12'sd1077, 12'sd-2026}},
{{12'sd1107, 12'sd-1136, 13'sd3909}, {13'sd3279, 12'sd-1680, 13'sd2050}, {14'sd4353, 12'sd-1253, 13'sd3810}},
{{9'sd-143, 12'sd1506, 12'sd-1578}, {12'sd-1300, 13'sd-2239, 10'sd480}, {13'sd2292, 10'sd281, 12'sd1959}},
{{14'sd-8047, 13'sd-3004, 14'sd-5765}, {12'sd-1957, 10'sd-325, 13'sd-3919}, {9'sd-250, 12'sd-1635, 13'sd-3229}},
{{12'sd1245, 13'sd2504, 12'sd1171}, {13'sd2925, 10'sd-418, 12'sd-1871}, {12'sd-1087, 13'sd-2645, 11'sd631}},
{{7'sd60, 9'sd-187, 13'sd3039}, {11'sd-622, 12'sd1194, 10'sd331}, {6'sd-22, 13'sd-2362, 13'sd2665}},
{{11'sd-578, 12'sd1155, 13'sd2591}, {13'sd-2478, 11'sd-711, 12'sd-1905}, {12'sd1303, 10'sd-390, 10'sd-502}},
{{7'sd51, 10'sd-451, 11'sd863}, {13'sd-2691, 8'sd80, 13'sd2189}, {12'sd-1800, 12'sd-1041, 9'sd252}},
{{6'sd-20, 9'sd-136, 9'sd183}, {11'sd692, 12'sd1872, 11'sd-980}, {9'sd216, 13'sd-2400, 11'sd583}},
{{12'sd-1998, 12'sd-1351, 10'sd-449}, {9'sd-215, 11'sd-993, 10'sd269}, {11'sd815, 10'sd-266, 9'sd-220}},
{{12'sd-1233, 10'sd498, 13'sd2787}, {13'sd3000, 13'sd3253, 13'sd3462}, {13'sd2738, 13'sd2356, 11'sd632}},
{{13'sd2437, 10'sd410, 12'sd-1109}, {13'sd-2274, 13'sd-2394, 12'sd-1446}, {11'sd-887, 11'sd630, 11'sd-983}},
{{12'sd-2009, 9'sd-188, 11'sd-750}, {12'sd1774, 11'sd582, 11'sd-544}, {6'sd22, 12'sd1154, 11'sd-663}},
{{12'sd-1822, 7'sd58, 11'sd-847}, {11'sd-832, 12'sd1658, 12'sd-1772}, {12'sd-1887, 12'sd-1141, 12'sd1577}},
{{13'sd-2192, 13'sd2630, 12'sd1852}, {12'sd1447, 10'sd-483, 12'sd1182}, {13'sd-3247, 11'sd798, 12'sd-1603}},
{{11'sd-816, 11'sd609, 12'sd1298}, {13'sd-2245, 10'sd-494, 12'sd1881}, {12'sd-1840, 12'sd-1261, 13'sd-3127}},
{{13'sd2059, 12'sd-1834, 13'sd-2058}, {13'sd-2118, 13'sd-2102, 13'sd-3451}, {13'sd3705, 13'sd3647, 12'sd1281}},
{{12'sd-1569, 12'sd1432, 10'sd443}, {10'sd296, 13'sd-2081, 5'sd12}, {12'sd1211, 12'sd1214, 13'sd-3281}},
{{12'sd-1185, 13'sd2521, 13'sd2769}, {13'sd2121, 12'sd-1032, 12'sd-1789}, {13'sd2345, 13'sd-2285, 11'sd-773}},
{{14'sd-4107, 13'sd-3495, 11'sd-589}, {10'sd-380, 10'sd-324, 12'sd1418}, {12'sd1179, 9'sd-198, 11'sd998}},
{{12'sd1199, 12'sd1207, 13'sd-2098}, {11'sd-952, 9'sd232, 11'sd-616}, {12'sd1508, 12'sd-1593, 12'sd-1819}},
{{13'sd-3752, 13'sd-2100, 12'sd1739}, {12'sd-1041, 11'sd-760, 12'sd-1358}, {13'sd-3170, 12'sd-1180, 12'sd-2015}},
{{11'sd-938, 11'sd534, 12'sd-1519}, {11'sd821, 11'sd-590, 12'sd-1630}, {13'sd-3570, 10'sd-264, 12'sd1814}},
{{13'sd2405, 13'sd-3279, 13'sd3470}, {14'sd5085, 11'sd-1000, 12'sd1111}, {10'sd361, 10'sd485, 8'sd-92}},
{{12'sd-1033, 12'sd-1189, 11'sd-800}, {12'sd-1288, 13'sd-2884, 11'sd-844}, {12'sd-1857, 11'sd-534, 11'sd-628}},
{{13'sd-2353, 12'sd-1232, 8'sd88}, {12'sd1572, 11'sd-921, 11'sd-524}, {11'sd658, 12'sd-1531, 12'sd2023}},
{{10'sd452, 12'sd-1033, 4'sd-4}, {10'sd-498, 11'sd885, 11'sd771}, {12'sd1703, 13'sd-2162, 13'sd-2231}},
{{12'sd-1774, 12'sd-1290, 13'sd-2947}, {11'sd-584, 13'sd-2458, 11'sd-760}, {9'sd-145, 12'sd1131, 11'sd922}},
{{13'sd2409, 11'sd546, 12'sd1886}, {13'sd3077, 12'sd1414, 12'sd-1903}, {12'sd-1869, 13'sd-2305, 9'sd253}},
{{9'sd-211, 12'sd-1286, 13'sd-2679}, {11'sd593, 12'sd-1622, 12'sd-1668}, {11'sd845, 8'sd-120, 13'sd-2253}},
{{13'sd-2763, 13'sd-2379, 12'sd-1189}, {12'sd1300, 11'sd-958, 10'sd496}, {13'sd3119, 12'sd1169, 13'sd2479}},
{{12'sd-2018, 13'sd-2795, 14'sd-4658}, {12'sd-1076, 10'sd-393, 13'sd-2850}, {12'sd2028, 13'sd2498, 12'sd-1633}},
{{8'sd74, 10'sd-313, 10'sd291}, {10'sd298, 13'sd-3062, 12'sd1599}, {11'sd839, 13'sd-3261, 9'sd166}},
{{13'sd-2325, 13'sd-2555, 13'sd3834}, {11'sd-615, 11'sd822, 10'sd477}, {8'sd107, 12'sd1960, 11'sd648}},
{{13'sd-2353, 9'sd146, 10'sd336}, {11'sd984, 13'sd3371, 10'sd490}, {12'sd1328, 12'sd1533, 11'sd-754}},
{{8'sd105, 11'sd-772, 11'sd965}, {13'sd2243, 12'sd2015, 11'sd556}, {11'sd-1002, 12'sd1108, 13'sd-2421}},
{{7'sd43, 10'sd-386, 10'sd-258}, {12'sd1076, 12'sd-1179, 12'sd-1684}, {10'sd-472, 13'sd2241, 13'sd-3005}},
{{12'sd-1813, 11'sd740, 12'sd-2019}, {11'sd-860, 13'sd-2662, 13'sd-3163}, {14'sd-7189, 12'sd-1114, 13'sd-3338}},
{{12'sd2002, 11'sd540, 9'sd-214}, {11'sd933, 13'sd-2208, 12'sd-1589}, {12'sd1984, 13'sd-2791, 13'sd2355}},
{{12'sd-1208, 12'sd-1132, 12'sd-1571}, {13'sd-3975, 12'sd-1222, 12'sd-1099}, {13'sd-2595, 12'sd-1318, 11'sd536}},
{{13'sd3293, 12'sd1355, 12'sd1830}, {10'sd-505, 10'sd-298, 12'sd-1738}, {13'sd2241, 13'sd3658, 13'sd2829}},
{{13'sd-2290, 13'sd-2323, 13'sd-2902}, {12'sd-1115, 12'sd2019, 12'sd-1175}, {11'sd-705, 12'sd-1356, 11'sd605}},
{{12'sd-1904, 13'sd-2048, 13'sd-2083}, {9'sd-130, 10'sd-465, 13'sd-3407}, {12'sd-1708, 12'sd-1542, 13'sd-3498}},
{{11'sd849, 12'sd-1418, 13'sd3222}, {13'sd2455, 9'sd-250, 12'sd-1460}, {12'sd-1375, 10'sd-366, 14'sd4328}},
{{13'sd2227, 11'sd876, 12'sd-1292}, {10'sd-342, 10'sd-509, 12'sd1681}, {9'sd251, 13'sd2956, 13'sd2335}},
{{13'sd-2539, 13'sd-2710, 14'sd-4406}, {14'sd-4196, 8'sd118, 13'sd-4092}, {13'sd-3849, 12'sd-1957, 12'sd-1683}},
{{8'sd108, 12'sd1535, 13'sd3297}, {11'sd-916, 13'sd-2249, 12'sd-1307}, {8'sd-68, 11'sd-890, 12'sd-1111}}},
{
{{13'sd2849, 12'sd1191, 11'sd-1013}, {12'sd-1600, 8'sd-70, 11'sd-655}, {13'sd2901, 11'sd-940, 11'sd753}},
{{12'sd1403, 12'sd-1609, 12'sd-1529}, {12'sd1871, 11'sd518, 7'sd40}, {12'sd-1024, 11'sd-521, 13'sd-2613}},
{{11'sd-1013, 13'sd3431, 13'sd3428}, {9'sd160, 11'sd-697, 13'sd2260}, {13'sd-2406, 13'sd-2985, 13'sd-3995}},
{{8'sd-73, 13'sd-2875, 13'sd-2621}, {13'sd-2129, 9'sd-199, 11'sd842}, {12'sd1291, 12'sd-1294, 13'sd2221}},
{{13'sd-2463, 11'sd513, 11'sd-701}, {13'sd2293, 10'sd376, 13'sd-2611}, {12'sd-1676, 13'sd2303, 12'sd-1800}},
{{12'sd1900, 13'sd-2050, 8'sd93}, {12'sd1303, 12'sd1661, 11'sd762}, {12'sd-1179, 11'sd-900, 13'sd-2583}},
{{12'sd1928, 13'sd-3560, 13'sd-2611}, {12'sd-1197, 11'sd-861, 12'sd1431}, {13'sd3453, 13'sd3169, 9'sd-152}},
{{12'sd-1943, 12'sd-1150, 13'sd-3139}, {11'sd-968, 12'sd1351, 12'sd-1554}, {11'sd-791, 12'sd1163, 12'sd-1713}},
{{13'sd-2623, 10'sd372, 12'sd1353}, {12'sd-1408, 12'sd-1553, 10'sd263}, {12'sd-1518, 13'sd-2710, 12'sd1377}},
{{11'sd-679, 12'sd1233, 11'sd607}, {10'sd-445, 13'sd-2572, 13'sd-2086}, {12'sd-1713, 12'sd-1407, 9'sd235}},
{{12'sd-1628, 12'sd-1405, 5'sd15}, {11'sd718, 12'sd1705, 12'sd1895}, {12'sd-1913, 11'sd-1023, 12'sd-1831}},
{{10'sd-308, 13'sd-2555, 11'sd832}, {9'sd-172, 11'sd588, 13'sd-2461}, {11'sd629, 13'sd-2359, 13'sd-2484}},
{{12'sd1908, 10'sd-337, 13'sd-2989}, {13'sd-2622, 11'sd-729, 13'sd-3824}, {11'sd632, 12'sd-1096, 13'sd-2271}},
{{12'sd1205, 10'sd387, 11'sd-610}, {9'sd242, 9'sd148, 9'sd213}, {11'sd-520, 12'sd-1914, 12'sd-1031}},
{{12'sd-2008, 13'sd-2942, 12'sd1982}, {12'sd1808, 10'sd-417, 7'sd-56}, {13'sd-2048, 13'sd-3070, 12'sd1315}},
{{12'sd1324, 9'sd-225, 11'sd718}, {13'sd-2625, 11'sd697, 13'sd2305}, {13'sd-2290, 9'sd227, 12'sd-1348}},
{{12'sd-1631, 12'sd-1260, 12'sd1157}, {11'sd642, 12'sd1340, 10'sd-332}, {13'sd-2632, 13'sd2523, 13'sd2124}},
{{10'sd414, 10'sd-306, 12'sd1186}, {11'sd-636, 7'sd55, 12'sd-1546}, {13'sd-2498, 12'sd1034, 10'sd-308}},
{{13'sd-3410, 10'sd-285, 13'sd-2062}, {10'sd-341, 10'sd-466, 7'sd-38}, {11'sd-684, 13'sd-2881, 12'sd1199}},
{{12'sd-1483, 12'sd-1779, 12'sd-1752}, {13'sd-2262, 12'sd-1970, 11'sd533}, {12'sd1485, 11'sd538, 12'sd-1605}},
{{8'sd70, 13'sd2411, 12'sd-1246}, {13'sd2828, 13'sd-2829, 12'sd-1932}, {9'sd-164, 2'sd-1, 13'sd2697}},
{{13'sd-2357, 11'sd596, 12'sd-1731}, {13'sd2429, 12'sd1591, 10'sd486}, {11'sd-785, 12'sd-1094, 12'sd1501}},
{{13'sd2166, 12'sd1617, 12'sd1961}, {11'sd953, 13'sd-2143, 12'sd-1665}, {12'sd1749, 11'sd-541, 12'sd-1502}},
{{13'sd-2386, 12'sd1954, 12'sd-2022}, {13'sd2828, 13'sd2065, 7'sd-57}, {13'sd2467, 10'sd298, 12'sd-1955}},
{{13'sd-2751, 9'sd-145, 9'sd225}, {12'sd1197, 10'sd477, 10'sd-433}, {8'sd-81, 12'sd-1361, 8'sd72}},
{{11'sd529, 12'sd1769, 13'sd-2146}, {13'sd2465, 12'sd1525, 12'sd-1697}, {12'sd-1134, 11'sd791, 11'sd950}},
{{11'sd736, 11'sd-871, 12'sd-1201}, {11'sd655, 12'sd1629, 10'sd335}, {9'sd-136, 13'sd-3014, 13'sd-2569}},
{{12'sd-1646, 11'sd-720, 12'sd-1473}, {13'sd-2893, 11'sd-631, 12'sd-1415}, {12'sd1139, 12'sd1363, 11'sd667}},
{{13'sd2463, 12'sd1367, 12'sd-1339}, {12'sd1379, 13'sd-2450, 9'sd224}, {13'sd-2110, 13'sd-2225, 12'sd-1979}},
{{12'sd-1476, 12'sd1205, 11'sd-848}, {12'sd-2036, 13'sd2510, 10'sd-385}, {12'sd1718, 13'sd2530, 12'sd1994}},
{{10'sd331, 12'sd1442, 10'sd-397}, {11'sd-861, 14'sd5173, 13'sd3217}, {13'sd-3093, 8'sd101, 11'sd624}},
{{11'sd-586, 11'sd993, 12'sd1236}, {12'sd1462, 11'sd999, 9'sd134}, {12'sd1486, 12'sd-1966, 10'sd-500}},
{{13'sd-2782, 12'sd-1413, 9'sd240}, {13'sd2460, 12'sd-1844, 12'sd-1118}, {6'sd23, 12'sd1809, 13'sd2887}},
{{12'sd1625, 12'sd-1110, 13'sd2984}, {12'sd1475, 7'sd-54, 12'sd-1248}, {10'sd-299, 12'sd-1029, 12'sd1052}},
{{12'sd1772, 12'sd-1059, 10'sd455}, {12'sd-1292, 8'sd-102, 11'sd-896}, {13'sd2832, 12'sd-1263, 11'sd-935}},
{{11'sd989, 13'sd2629, 11'sd-525}, {7'sd-60, 11'sd-592, 6'sd16}, {12'sd-1596, 13'sd-2426, 12'sd1499}},
{{12'sd-1650, 9'sd192, 13'sd2279}, {11'sd998, 9'sd-175, 9'sd-195}, {11'sd-988, 12'sd1090, 12'sd1785}},
{{12'sd1575, 12'sd-1562, 9'sd-204}, {9'sd-197, 7'sd-36, 11'sd-844}, {11'sd769, 11'sd641, 12'sd-1222}},
{{11'sd-514, 12'sd-1585, 10'sd455}, {9'sd201, 7'sd38, 11'sd-733}, {11'sd-642, 13'sd2060, 12'sd-1786}},
{{13'sd-2422, 12'sd1419, 11'sd-1016}, {11'sd-993, 11'sd-1016, 11'sd952}, {12'sd1468, 12'sd1313, 12'sd1507}},
{{13'sd-3867, 12'sd1564, 10'sd309}, {12'sd1344, 11'sd-943, 12'sd1099}, {14'sd4114, 14'sd4204, 13'sd3377}},
{{13'sd2801, 13'sd3237, 12'sd1658}, {13'sd2082, 12'sd1411, 12'sd-1700}, {6'sd27, 9'sd249, 12'sd-1740}},
{{12'sd-1473, 13'sd-2183, 9'sd-176}, {10'sd-367, 12'sd-2007, 11'sd522}, {13'sd3316, 11'sd649, 11'sd698}},
{{13'sd-2701, 11'sd912, 12'sd-1222}, {13'sd2153, 12'sd1792, 12'sd1710}, {12'sd1280, 10'sd395, 13'sd-2075}},
{{11'sd-608, 7'sd-47, 8'sd72}, {12'sd-1650, 13'sd2196, 9'sd-138}, {8'sd72, 11'sd-540, 13'sd-2191}},
{{13'sd-2712, 12'sd-1426, 10'sd275}, {9'sd-238, 12'sd-1932, 12'sd1948}, {13'sd2416, 13'sd2163, 12'sd-1709}},
{{10'sd317, 13'sd-2216, 11'sd-737}, {8'sd93, 12'sd-1627, 12'sd-1481}, {13'sd2059, 12'sd2017, 9'sd149}},
{{14'sd4141, 13'sd3520, 12'sd1626}, {12'sd1653, 10'sd-256, 11'sd-947}, {12'sd-1528, 12'sd1232, 13'sd2457}},
{{12'sd1590, 14'sd4699, 12'sd1661}, {13'sd-2752, 13'sd2805, 11'sd-982}, {12'sd-1999, 13'sd3891, 13'sd2083}},
{{13'sd-3416, 13'sd-2396, 11'sd-757}, {8'sd-113, 12'sd-1452, 12'sd-1403}, {12'sd-1758, 13'sd2624, 12'sd1277}},
{{13'sd2734, 13'sd2056, 12'sd-1785}, {13'sd2793, 11'sd834, 13'sd2494}, {11'sd887, 11'sd567, 13'sd-2351}},
{{13'sd2142, 11'sd701, 13'sd-2539}, {12'sd1170, 11'sd-948, 12'sd1465}, {11'sd-767, 13'sd-2922, 11'sd562}},
{{8'sd85, 13'sd-2606, 13'sd-2626}, {13'sd2501, 11'sd946, 13'sd2680}, {11'sd551, 10'sd-421, 12'sd-1703}},
{{12'sd1791, 13'sd2193, 13'sd-2466}, {12'sd-2007, 11'sd-892, 11'sd737}, {11'sd-663, 9'sd-171, 12'sd-1820}},
{{14'sd5440, 13'sd3897, 8'sd-97}, {13'sd3720, 12'sd1344, 13'sd-2301}, {9'sd-156, 12'sd-1754, 13'sd-3525}},
{{10'sd-441, 9'sd163, 11'sd601}, {10'sd-269, 12'sd1971, 12'sd-1658}, {13'sd2167, 11'sd788, 12'sd-1270}},
{{10'sd-479, 12'sd1223, 12'sd1847}, {12'sd2042, 13'sd2604, 11'sd700}, {12'sd1128, 12'sd1114, 13'sd-2436}},
{{12'sd1823, 13'sd-2278, 13'sd2570}, {13'sd-2072, 11'sd-632, 12'sd1146}, {11'sd-843, 13'sd-3221, 11'sd-651}},
{{11'sd760, 12'sd-1802, 11'sd-897}, {13'sd2687, 12'sd1541, 13'sd-2343}, {13'sd2329, 10'sd415, 13'sd3359}},
{{14'sd4146, 13'sd2266, 12'sd1917}, {12'sd1401, 12'sd1400, 10'sd291}, {12'sd-1762, 12'sd1179, 10'sd-369}},
{{11'sd982, 12'sd1205, 12'sd1203}, {10'sd391, 12'sd1039, 12'sd1273}, {10'sd349, 12'sd-1066, 12'sd1825}},
{{6'sd-23, 12'sd1639, 11'sd-545}, {13'sd-2918, 13'sd3620, 13'sd2430}, {10'sd352, 9'sd155, 11'sd821}},
{{13'sd3360, 13'sd2152, 13'sd3250}, {13'sd2548, 12'sd-1444, 12'sd1181}, {12'sd1096, 13'sd-2296, 12'sd1248}},
{{12'sd1224, 12'sd1152, 11'sd643}, {12'sd-1734, 13'sd3366, 4'sd-7}, {12'sd-1051, 11'sd844, 12'sd1928}}},
{
{{12'sd1456, 13'sd-2445, 13'sd-2438}, {12'sd1029, 11'sd-786, 13'sd-2228}, {13'sd2261, 12'sd-1559, 10'sd-411}},
{{13'sd2696, 12'sd1689, 5'sd-8}, {13'sd-2161, 11'sd942, 12'sd-1344}, {10'sd-278, 12'sd-1160, 12'sd1976}},
{{11'sd-959, 11'sd-825, 10'sd-377}, {12'sd1310, 10'sd-339, 11'sd-681}, {11'sd938, 13'sd2702, 13'sd2630}},
{{9'sd-203, 12'sd-1723, 11'sd559}, {10'sd510, 12'sd-1824, 12'sd-1556}, {12'sd1489, 10'sd383, 12'sd1233}},
{{12'sd1277, 10'sd407, 9'sd-235}, {10'sd-439, 13'sd-2325, 12'sd-1525}, {13'sd-2443, 12'sd-1266, 11'sd-666}},
{{12'sd1719, 10'sd485, 12'sd-1465}, {11'sd-706, 11'sd1006, 13'sd-2366}, {13'sd2212, 12'sd-1802, 8'sd73}},
{{9'sd168, 10'sd-303, 12'sd-2001}, {13'sd2784, 8'sd-85, 13'sd-2212}, {13'sd-2155, 13'sd-2749, 12'sd-1216}},
{{11'sd678, 11'sd590, 12'sd-1493}, {13'sd-2237, 12'sd1984, 12'sd1075}, {11'sd-915, 13'sd2441, 10'sd336}},
{{13'sd-2127, 12'sd1049, 11'sd-686}, {12'sd1891, 10'sd491, 10'sd-378}, {11'sd-594, 12'sd-1999, 10'sd491}},
{{12'sd1843, 12'sd-1812, 11'sd-588}, {11'sd-529, 8'sd-113, 10'sd-345}, {9'sd-230, 12'sd-1152, 12'sd-1383}},
{{13'sd-2235, 12'sd1368, 11'sd656}, {11'sd839, 9'sd217, 12'sd1716}, {13'sd2676, 9'sd184, 11'sd-907}},
{{13'sd2596, 12'sd1922, 13'sd2713}, {12'sd-1775, 13'sd-2268, 13'sd2177}, {12'sd1134, 11'sd580, 12'sd1725}},
{{9'sd-227, 13'sd3591, 11'sd-945}, {10'sd-352, 11'sd804, 13'sd-2615}, {12'sd2013, 13'sd-3573, 11'sd-983}},
{{12'sd1699, 11'sd1018, 12'sd1922}, {11'sd-683, 13'sd2300, 13'sd-2148}, {11'sd-880, 13'sd-2754, 12'sd1119}},
{{12'sd-1266, 12'sd1662, 11'sd756}, {12'sd-1652, 10'sd-449, 13'sd-2138}, {13'sd2647, 9'sd-193, 12'sd-1194}},
{{11'sd762, 8'sd-115, 13'sd2793}, {13'sd2234, 12'sd1742, 12'sd1958}, {11'sd859, 12'sd1857, 11'sd630}},
{{13'sd-2609, 13'sd2366, 13'sd2740}, {10'sd383, 10'sd-487, 12'sd1592}, {10'sd262, 12'sd1039, 9'sd182}},
{{14'sd-4831, 13'sd-3064, 11'sd603}, {12'sd1228, 11'sd-808, 13'sd2314}, {13'sd-2365, 13'sd2774, 13'sd2980}},
{{12'sd1276, 12'sd-1725, 13'sd2095}, {12'sd-1061, 13'sd2567, 13'sd-2910}, {12'sd-1450, 12'sd-1356, 11'sd-801}},
{{12'sd1517, 13'sd2687, 11'sd-1017}, {11'sd-574, 12'sd1522, 12'sd1265}, {11'sd866, 11'sd885, 12'sd-1948}},
{{12'sd-1281, 13'sd2472, 12'sd-1791}, {13'sd-2263, 12'sd-1550, 12'sd-1411}, {13'sd2343, 12'sd1181, 12'sd-1324}},
{{13'sd-2737, 13'sd2347, 12'sd1450}, {12'sd-1770, 11'sd948, 12'sd1997}, {12'sd1857, 12'sd-1905, 11'sd720}},
{{9'sd-205, 12'sd-1261, 12'sd1329}, {12'sd1296, 12'sd-1383, 13'sd-2156}, {12'sd1134, 13'sd2402, 8'sd105}},
{{12'sd-1829, 13'sd-2333, 12'sd1252}, {9'sd-176, 12'sd1746, 12'sd1165}, {11'sd588, 12'sd-1874, 11'sd804}},
{{10'sd355, 11'sd600, 11'sd-911}, {12'sd1127, 10'sd-282, 10'sd495}, {11'sd-782, 12'sd1509, 12'sd2034}},
{{13'sd2487, 10'sd-452, 12'sd-1783}, {13'sd2649, 12'sd1723, 12'sd1841}, {13'sd2248, 12'sd1345, 11'sd682}},
{{9'sd164, 13'sd-2789, 12'sd1694}, {13'sd-3056, 10'sd-357, 11'sd-770}, {11'sd-917, 12'sd1376, 13'sd-2626}},
{{13'sd2592, 12'sd-1368, 13'sd-3147}, {10'sd327, 13'sd2328, 12'sd-1298}, {11'sd837, 12'sd1759, 13'sd-2725}},
{{13'sd2888, 11'sd-1023, 13'sd2606}, {13'sd2976, 12'sd-1794, 4'sd-5}, {10'sd-425, 12'sd1401, 13'sd2442}},
{{12'sd-1254, 13'sd-2055, 12'sd-1175}, {12'sd1923, 13'sd2666, 13'sd2347}, {12'sd-1847, 12'sd1426, 13'sd-2222}},
{{13'sd-3858, 9'sd201, 12'sd-1519}, {12'sd-1109, 12'sd-1659, 13'sd2529}, {14'sd-4714, 11'sd-518, 11'sd-589}},
{{12'sd1168, 11'sd-968, 13'sd-2251}, {12'sd-1927, 12'sd1947, 12'sd1055}, {9'sd-208, 11'sd-542, 12'sd1711}},
{{13'sd-3419, 11'sd-709, 12'sd-1823}, {12'sd-1366, 13'sd-3029, 10'sd-484}, {13'sd-3797, 13'sd-3842, 12'sd1861}},
{{12'sd-1535, 11'sd846, 13'sd2583}, {12'sd1696, 12'sd-1768, 12'sd1248}, {9'sd231, 12'sd2008, 13'sd2839}},
{{8'sd78, 9'sd-212, 12'sd1856}, {12'sd-1491, 10'sd-401, 12'sd-1413}, {11'sd-822, 13'sd2365, 12'sd-1836}},
{{12'sd1099, 13'sd2184, 12'sd-1901}, {12'sd-1921, 11'sd-542, 11'sd1020}, {10'sd322, 12'sd1057, 11'sd-864}},
{{12'sd-1761, 12'sd-2001, 11'sd1005}, {11'sd-963, 11'sd758, 9'sd-255}, {13'sd-2479, 11'sd-836, 12'sd-1405}},
{{11'sd-851, 12'sd1942, 7'sd45}, {11'sd-790, 13'sd-2436, 12'sd1711}, {13'sd2048, 13'sd-2319, 13'sd-2101}},
{{13'sd2258, 12'sd1339, 13'sd2256}, {12'sd1986, 10'sd-388, 13'sd-2266}, {11'sd989, 8'sd90, 13'sd-2202}},
{{12'sd1802, 13'sd-2957, 13'sd-2575}, {12'sd1822, 13'sd-2933, 12'sd-1604}, {11'sd-740, 13'sd-2170, 13'sd-2702}},
{{12'sd1957, 12'sd-1464, 13'sd-2089}, {13'sd2401, 10'sd474, 12'sd-2026}, {13'sd-2318, 12'sd1244, 13'sd-2726}},
{{13'sd3159, 13'sd3305, 12'sd-1464}, {12'sd1251, 12'sd1140, 9'sd-255}, {12'sd-1620, 11'sd-1009, 12'sd1598}},
{{10'sd-324, 12'sd1631, 11'sd606}, {8'sd-127, 12'sd-1392, 12'sd1843}, {12'sd1041, 13'sd2655, 5'sd-15}},
{{12'sd1952, 13'sd2162, 12'sd1085}, {11'sd-642, 12'sd1148, 13'sd2171}, {10'sd333, 13'sd2587, 12'sd-1533}},
{{10'sd457, 12'sd1195, 13'sd2580}, {13'sd2762, 11'sd-769, 12'sd-1806}, {13'sd3418, 12'sd-1907, 8'sd116}},
{{6'sd-22, 10'sd361, 9'sd-139}, {10'sd342, 11'sd789, 12'sd-1045}, {13'sd-2284, 13'sd3085, 10'sd-434}},
{{9'sd216, 11'sd-998, 12'sd-1142}, {13'sd2479, 11'sd534, 13'sd3033}, {12'sd-1269, 13'sd2903, 12'sd1890}},
{{12'sd1658, 11'sd512, 13'sd2710}, {12'sd-1396, 12'sd-1923, 12'sd-1664}, {12'sd1551, 12'sd1670, 8'sd82}},
{{13'sd-2096, 10'sd-411, 13'sd3076}, {13'sd-2220, 9'sd163, 11'sd-536}, {11'sd885, 10'sd328, 9'sd191}},
{{13'sd-2870, 11'sd614, 12'sd-1329}, {10'sd-293, 1'sd0, 13'sd2129}, {9'sd-213, 13'sd2198, 11'sd-701}},
{{14'sd4237, 12'sd1615, 13'sd-3313}, {9'sd-149, 13'sd-2511, 12'sd1087}, {12'sd-1533, 11'sd-692, 11'sd988}},
{{12'sd1728, 12'sd-1760, 12'sd-1529}, {13'sd-2431, 13'sd-2244, 11'sd802}, {12'sd1882, 12'sd-1790, 10'sd-500}},
{{13'sd-2591, 11'sd-634, 10'sd282}, {11'sd-643, 13'sd-2326, 12'sd1030}, {12'sd1196, 13'sd2591, 9'sd-230}},
{{12'sd-1456, 12'sd-1819, 12'sd-1668}, {11'sd-817, 11'sd-722, 13'sd-2350}, {11'sd727, 12'sd1038, 13'sd2121}},
{{12'sd1368, 13'sd2077, 10'sd388}, {9'sd-204, 10'sd-280, 12'sd1274}, {10'sd390, 13'sd-2616, 13'sd2278}},
{{13'sd2071, 11'sd-602, 11'sd621}, {12'sd1971, 13'sd3029, 11'sd568}, {11'sd-607, 12'sd1071, 11'sd686}},
{{12'sd-1925, 12'sd-1673, 9'sd186}, {11'sd709, 12'sd-1527, 11'sd-660}, {11'sd679, 11'sd702, 12'sd1573}},
{{9'sd-204, 12'sd1190, 11'sd574}, {11'sd-605, 12'sd-1041, 11'sd-746}, {13'sd2547, 13'sd2327, 8'sd-94}},
{{12'sd-2038, 11'sd-637, 12'sd-1908}, {12'sd-1770, 13'sd2200, 13'sd-2228}, {13'sd-3148, 13'sd-2866, 12'sd1503}},
{{13'sd3131, 13'sd3202, 12'sd-1194}, {11'sd817, 12'sd-1582, 11'sd952}, {7'sd-45, 12'sd-1146, 12'sd1074}},
{{12'sd1097, 4'sd6, 12'sd1133}, {12'sd1049, 12'sd-1157, 12'sd1301}, {9'sd-236, 11'sd-868, 9'sd-250}},
{{13'sd-2630, 8'sd77, 13'sd2122}, {12'sd-1058, 7'sd39, 12'sd1121}, {13'sd-2546, 11'sd828, 12'sd-1150}},
{{12'sd1729, 13'sd2328, 12'sd-1663}, {12'sd1241, 12'sd1115, 11'sd814}, {11'sd-710, 11'sd900, 13'sd-2229}},
{{6'sd22, 13'sd-2188, 12'sd-1839}, {11'sd621, 8'sd-106, 9'sd-239}, {6'sd25, 9'sd-190, 13'sd3001}}},
{
{{12'sd-1820, 10'sd-397, 8'sd-106}, {13'sd3100, 13'sd-2177, 13'sd2555}, {12'sd1224, 8'sd101, 13'sd3692}},
{{13'sd2614, 12'sd1833, 12'sd1737}, {8'sd-65, 11'sd-808, 11'sd762}, {13'sd2486, 11'sd531, 12'sd-1736}},
{{12'sd-1435, 12'sd-1888, 13'sd-2536}, {12'sd-1346, 10'sd497, 12'sd-1249}, {13'sd2352, 13'sd-2843, 12'sd1152}},
{{12'sd2040, 12'sd-1245, 13'sd2605}, {12'sd-1375, 12'sd1565, 12'sd-1303}, {12'sd-1659, 12'sd-1940, 13'sd2316}},
{{6'sd-31, 13'sd-2568, 13'sd2630}, {13'sd-3035, 13'sd-2393, 13'sd-2669}, {12'sd-1870, 10'sd-429, 12'sd1105}},
{{10'sd390, 12'sd1637, 13'sd-2132}, {12'sd-1254, 12'sd1814, 12'sd-1570}, {13'sd2351, 7'sd-43, 12'sd1668}},
{{12'sd1935, 12'sd-1618, 10'sd464}, {11'sd-885, 12'sd-1157, 12'sd1466}, {13'sd-3694, 12'sd-1809, 13'sd2672}},
{{12'sd-1929, 13'sd-2306, 12'sd-1820}, {10'sd-480, 12'sd-1785, 11'sd-523}, {12'sd2015, 13'sd-3034, 12'sd-1632}},
{{13'sd2202, 13'sd-2648, 11'sd891}, {12'sd1566, 10'sd-445, 12'sd2036}, {12'sd-1894, 12'sd1956, 10'sd502}},
{{13'sd-2426, 12'sd-1795, 12'sd-1691}, {12'sd1377, 10'sd-355, 12'sd-1558}, {12'sd-2023, 7'sd-48, 13'sd-2377}},
{{11'sd-593, 10'sd465, 12'sd1754}, {13'sd-2065, 12'sd-1400, 12'sd1568}, {13'sd2813, 13'sd2793, 13'sd2231}},
{{13'sd3587, 11'sd994, 12'sd-1595}, {12'sd-1981, 13'sd2803, 11'sd-817}, {13'sd3184, 12'sd1680, 10'sd493}},
{{13'sd3063, 12'sd1069, 13'sd3965}, {13'sd2831, 13'sd2472, 11'sd-858}, {12'sd-1491, 13'sd2627, 12'sd-1972}},
{{11'sd686, 13'sd2592, 10'sd-445}, {13'sd2250, 12'sd2029, 11'sd752}, {12'sd-1773, 12'sd-1291, 13'sd3015}},
{{12'sd-1123, 8'sd-114, 13'sd-2867}, {13'sd2306, 12'sd1093, 13'sd2365}, {13'sd-2597, 11'sd805, 12'sd1232}},
{{11'sd958, 11'sd871, 11'sd-918}, {13'sd-2425, 9'sd-182, 13'sd-2481}, {9'sd193, 12'sd-1386, 12'sd2009}},
{{11'sd-706, 11'sd-558, 11'sd-722}, {10'sd459, 12'sd-1247, 10'sd-375}, {12'sd1679, 13'sd2104, 9'sd153}},
{{11'sd-951, 10'sd508, 13'sd3382}, {13'sd-2524, 12'sd-1139, 12'sd1928}, {11'sd978, 12'sd-1614, 13'sd3861}},
{{9'sd-236, 9'sd236, 13'sd2334}, {12'sd1640, 11'sd930, 6'sd-24}, {11'sd928, 11'sd-864, 11'sd-964}},
{{12'sd1707, 12'sd-1413, 11'sd597}, {12'sd-1163, 10'sd374, 10'sd511}, {11'sd767, 12'sd-1338, 12'sd-1492}},
{{12'sd1566, 11'sd-826, 9'sd162}, {6'sd-21, 13'sd-2479, 11'sd949}, {12'sd-1945, 7'sd36, 13'sd2124}},
{{11'sd829, 13'sd2976, 12'sd-1996}, {12'sd1485, 13'sd2313, 9'sd185}, {9'sd230, 11'sd-809, 12'sd-1294}},
{{11'sd555, 12'sd1312, 13'sd2301}, {12'sd-1395, 12'sd-1057, 12'sd1703}, {12'sd1935, 12'sd1115, 13'sd2217}},
{{12'sd-1705, 11'sd-688, 12'sd1418}, {9'sd-160, 12'sd-1997, 13'sd-2171}, {13'sd-2600, 13'sd-3327, 8'sd108}},
{{12'sd-1103, 13'sd2119, 12'sd-1146}, {8'sd-98, 13'sd2063, 9'sd-232}, {8'sd-110, 13'sd-2146, 13'sd2309}},
{{13'sd-2413, 10'sd-316, 12'sd1657}, {11'sd981, 12'sd1078, 7'sd50}, {13'sd2462, 10'sd-415, 12'sd-1792}},
{{12'sd-1117, 13'sd2187, 7'sd38}, {12'sd-1991, 11'sd-957, 13'sd-2393}, {11'sd-947, 11'sd669, 13'sd-2308}},
{{13'sd2521, 12'sd-1510, 10'sd371}, {8'sd82, 13'sd2346, 12'sd1407}, {13'sd-3534, 13'sd-2658, 11'sd564}},
{{12'sd-1819, 13'sd2209, 10'sd-316}, {10'sd-345, 12'sd-1771, 13'sd-2345}, {12'sd1275, 12'sd-1316, 11'sd897}},
{{12'sd1810, 12'sd-1543, 12'sd-1478}, {10'sd301, 13'sd2990, 11'sd748}, {11'sd784, 10'sd405, 13'sd-2831}},
{{13'sd-2802, 12'sd1919, 11'sd-712}, {13'sd-3261, 13'sd-2211, 9'sd217}, {13'sd-3047, 13'sd-2289, 11'sd-989}},
{{12'sd-1292, 10'sd507, 13'sd2304}, {11'sd620, 12'sd1542, 12'sd-1601}, {13'sd3029, 12'sd1551, 12'sd1922}},
{{7'sd-47, 13'sd2253, 12'sd-1484}, {11'sd998, 12'sd-2022, 13'sd4055}, {11'sd664, 13'sd-2680, 10'sd-327}},
{{12'sd1125, 12'sd-1451, 13'sd-3088}, {10'sd-407, 12'sd-1659, 12'sd-1347}, {13'sd-2826, 6'sd23, 13'sd-4067}},
{{13'sd-2455, 13'sd2100, 12'sd1263}, {12'sd1632, 12'sd1957, 11'sd-770}, {12'sd-1104, 13'sd2070, 13'sd2663}},
{{13'sd2789, 11'sd843, 12'sd1994}, {10'sd-418, 13'sd2092, 9'sd-220}, {11'sd-893, 4'sd-5, 11'sd-604}},
{{13'sd-2073, 11'sd-597, 10'sd-456}, {12'sd-1397, 11'sd548, 12'sd1031}, {12'sd1180, 10'sd489, 13'sd-2245}},
{{13'sd2586, 4'sd4, 13'sd-2506}, {12'sd-1227, 13'sd2554, 13'sd2191}, {12'sd1258, 13'sd2685, 13'sd-2350}},
{{12'sd1267, 10'sd469, 13'sd2340}, {12'sd1116, 11'sd-823, 10'sd502}, {10'sd-374, 13'sd2204, 9'sd-160}},
{{12'sd1262, 8'sd-66, 13'sd-2075}, {12'sd-1732, 12'sd-1361, 12'sd1858}, {12'sd-1546, 12'sd-1379, 12'sd-1324}},
{{14'sd4216, 12'sd-1243, 13'sd2556}, {11'sd768, 12'sd-2013, 13'sd3219}, {11'sd927, 13'sd2874, 14'sd4164}},
{{12'sd-1943, 12'sd1098, 11'sd-730}, {11'sd-885, 12'sd-1218, 12'sd1773}, {11'sd-850, 12'sd2000, 12'sd1616}},
{{11'sd795, 12'sd-1853, 12'sd1121}, {13'sd2511, 13'sd2839, 13'sd-2292}, {13'sd3460, 13'sd2459, 13'sd2633}},
{{12'sd-1843, 13'sd2888, 13'sd-2131}, {13'sd-2710, 11'sd799, 11'sd-709}, {11'sd692, 13'sd-2084, 11'sd850}},
{{11'sd546, 10'sd-446, 13'sd2284}, {13'sd2550, 5'sd-13, 11'sd-849}, {11'sd-810, 13'sd-2607, 13'sd-2559}},
{{12'sd-1354, 12'sd-1478, 13'sd2549}, {12'sd1699, 11'sd808, 13'sd2219}, {13'sd2472, 13'sd2940, 13'sd2062}},
{{13'sd2826, 11'sd-828, 10'sd486}, {13'sd2630, 11'sd-604, 11'sd961}, {12'sd1031, 12'sd1751, 13'sd2544}},
{{12'sd1569, 13'sd2410, 13'sd2396}, {13'sd2326, 8'sd71, 9'sd219}, {13'sd3202, 13'sd3399, 12'sd-1688}},
{{13'sd-3628, 13'sd2201, 13'sd2422}, {14'sd-4583, 13'sd-3028, 13'sd2251}, {13'sd-3673, 12'sd-1755, 11'sd-827}},
{{12'sd1900, 6'sd-25, 13'sd2506}, {12'sd-1730, 12'sd-1243, 12'sd1268}, {10'sd-421, 9'sd251, 11'sd-663}},
{{12'sd-1481, 12'sd-1058, 11'sd726}, {12'sd-1180, 12'sd2002, 13'sd-2401}, {12'sd1873, 12'sd-1405, 11'sd-585}},
{{12'sd-1842, 13'sd2928, 12'sd1330}, {12'sd-1931, 12'sd-1191, 13'sd2616}, {8'sd-69, 11'sd-767, 7'sd41}},
{{13'sd2579, 12'sd-1623, 13'sd-2586}, {10'sd-325, 10'sd-327, 13'sd-2956}, {12'sd1321, 11'sd-829, 13'sd-3139}},
{{11'sd-763, 11'sd978, 13'sd2653}, {13'sd-3049, 10'sd339, 11'sd-818}, {11'sd911, 10'sd434, 12'sd1432}},
{{12'sd1420, 13'sd3462, 13'sd-2392}, {11'sd-633, 10'sd-262, 11'sd593}, {13'sd2196, 9'sd-213, 12'sd1416}},
{{11'sd-741, 12'sd-2038, 12'sd-1774}, {12'sd1151, 12'sd-1773, 11'sd749}, {12'sd1714, 11'sd-593, 10'sd381}},
{{11'sd-525, 12'sd-1512, 13'sd2615}, {12'sd1851, 11'sd-632, 12'sd1050}, {11'sd761, 13'sd-2220, 11'sd-995}},
{{13'sd2403, 9'sd249, 11'sd836}, {11'sd-616, 13'sd2328, 12'sd1853}, {9'sd-227, 11'sd589, 13'sd-2288}},
{{12'sd-1306, 13'sd3030, 10'sd-328}, {12'sd1079, 13'sd-2055, 10'sd-399}, {12'sd1277, 12'sd1078, 12'sd1180}},
{{13'sd2415, 11'sd-803, 12'sd-1242}, {5'sd-15, 12'sd1190, 12'sd-1847}, {10'sd-299, 10'sd-496, 12'sd-1196}},
{{13'sd2920, 12'sd1073, 11'sd763}, {12'sd1399, 13'sd-2958, 12'sd1778}, {11'sd807, 8'sd-78, 12'sd-1698}},
{{12'sd-1291, 9'sd224, 12'sd-1168}, {11'sd-776, 8'sd-117, 9'sd-217}, {13'sd-2142, 13'sd-2557, 13'sd2532}},
{{11'sd927, 12'sd-1963, 9'sd-171}, {13'sd-2392, 13'sd-2515, 10'sd-337}, {11'sd910, 11'sd-695, 12'sd-1127}},
{{12'sd1239, 13'sd2254, 12'sd1663}, {12'sd1544, 11'sd943, 12'sd-1436}, {12'sd1458, 11'sd1013, 12'sd-1255}}},
{
{{13'sd-3106, 11'sd527, 6'sd-30}, {13'sd-2609, 11'sd-962, 13'sd-2399}, {13'sd-2077, 13'sd-2413, 10'sd383}},
{{12'sd-1047, 12'sd1685, 13'sd2463}, {12'sd1999, 13'sd2745, 9'sd158}, {13'sd-3221, 9'sd-142, 10'sd-355}},
{{10'sd-448, 11'sd-559, 12'sd-1783}, {12'sd-1588, 9'sd192, 12'sd1605}, {11'sd933, 11'sd772, 12'sd1580}},
{{11'sd-536, 12'sd1123, 12'sd1269}, {9'sd222, 10'sd-308, 11'sd-769}, {12'sd1792, 12'sd1530, 11'sd906}},
{{11'sd743, 12'sd-1186, 13'sd3271}, {11'sd-615, 12'sd-1270, 10'sd277}, {13'sd2329, 12'sd-1186, 12'sd1701}},
{{12'sd1317, 12'sd2015, 13'sd-2213}, {12'sd-1362, 12'sd-1226, 12'sd-1504}, {11'sd-863, 10'sd297, 11'sd567}},
{{12'sd-1691, 12'sd1071, 9'sd162}, {12'sd1104, 11'sd-719, 12'sd1203}, {11'sd878, 6'sd-21, 12'sd-1348}},
{{12'sd-1236, 13'sd-3448, 13'sd-2671}, {8'sd73, 12'sd-1394, 12'sd-1282}, {13'sd-2243, 11'sd-837, 12'sd1915}},
{{12'sd1166, 12'sd-1408, 9'sd-185}, {11'sd-906, 13'sd2232, 12'sd1127}, {12'sd-1359, 12'sd-1240, 12'sd1092}},
{{11'sd857, 12'sd1822, 10'sd346}, {9'sd255, 12'sd1977, 13'sd2321}, {13'sd2425, 12'sd2010, 11'sd-738}},
{{12'sd-1400, 5'sd-10, 11'sd-631}, {12'sd-1575, 12'sd1417, 12'sd1773}, {11'sd738, 10'sd285, 11'sd-742}},
{{10'sd-464, 8'sd66, 13'sd-3884}, {12'sd1246, 12'sd-1431, 12'sd1468}, {12'sd-1662, 11'sd1002, 12'sd-1926}},
{{13'sd-2982, 9'sd237, 11'sd968}, {12'sd1954, 11'sd-974, 12'sd1494}, {12'sd-1850, 11'sd-586, 11'sd947}},
{{12'sd2026, 8'sd-110, 12'sd1931}, {12'sd-1965, 12'sd-1911, 10'sd305}, {12'sd-1597, 12'sd1072, 12'sd1130}},
{{12'sd2024, 11'sd953, 13'sd-2908}, {12'sd-1461, 13'sd-2232, 10'sd450}, {7'sd32, 10'sd499, 13'sd-2137}},
{{13'sd3765, 10'sd465, 12'sd-1825}, {13'sd2953, 12'sd-1961, 12'sd-1492}, {13'sd3720, 12'sd1622, 9'sd-212}},
{{11'sd-560, 13'sd2119, 13'sd-2766}, {11'sd-520, 12'sd-2043, 12'sd1855}, {12'sd1230, 13'sd-3006, 13'sd-2883}},
{{13'sd3710, 11'sd643, 13'sd-2869}, {10'sd-266, 10'sd482, 13'sd-3115}, {14'sd4894, 13'sd3079, 13'sd2303}},
{{13'sd3349, 12'sd-1798, 11'sd-861}, {12'sd1761, 13'sd2996, 13'sd2162}, {12'sd1701, 13'sd2733, 10'sd-380}},
{{12'sd-1960, 13'sd2363, 13'sd2475}, {11'sd-645, 11'sd-850, 11'sd-664}, {10'sd281, 12'sd-1723, 13'sd2686}},
{{12'sd-1521, 11'sd-630, 12'sd1053}, {12'sd1316, 12'sd-1840, 13'sd2616}, {12'sd-1325, 13'sd-2635, 13'sd-3175}},
{{13'sd-3202, 11'sd615, 12'sd-1643}, {9'sd-202, 12'sd1197, 11'sd805}, {11'sd-564, 13'sd2743, 12'sd1062}},
{{12'sd1415, 8'sd-113, 10'sd-366}, {11'sd-822, 13'sd3111, 11'sd-713}, {13'sd2325, 12'sd-1894, 12'sd-1332}},
{{13'sd3149, 11'sd-746, 12'sd-1456}, {10'sd-261, 12'sd1058, 13'sd-2259}, {10'sd-263, 12'sd-1744, 9'sd-253}},
{{12'sd-1845, 13'sd-2088, 11'sd833}, {13'sd-2291, 13'sd-2880, 13'sd-2247}, {11'sd-762, 10'sd-343, 10'sd395}},
{{12'sd-1871, 11'sd-963, 11'sd-771}, {13'sd2561, 13'sd-2476, 13'sd2338}, {12'sd1665, 12'sd1996, 12'sd-1173}},
{{11'sd-621, 11'sd-772, 12'sd1821}, {13'sd2180, 11'sd673, 13'sd2435}, {12'sd1918, 11'sd986, 13'sd-2256}},
{{12'sd1810, 11'sd900, 14'sd4381}, {11'sd-804, 12'sd-1583, 12'sd-1466}, {10'sd420, 9'sd-238, 13'sd2601}},
{{11'sd-867, 7'sd33, 11'sd-926}, {12'sd1301, 10'sd-504, 12'sd1112}, {12'sd-1164, 12'sd1876, 13'sd2152}},
{{12'sd-1376, 13'sd3842, 13'sd2948}, {11'sd-891, 12'sd-2033, 12'sd-1110}, {12'sd2030, 10'sd300, 12'sd-1379}},
{{12'sd1815, 10'sd267, 11'sd-933}, {13'sd3896, 13'sd-2790, 13'sd-3824}, {14'sd4855, 12'sd1842, 13'sd-3686}},
{{13'sd-3074, 12'sd-1977, 13'sd-3192}, {13'sd-2780, 12'sd-1212, 8'sd83}, {12'sd-1046, 13'sd-2508, 11'sd-540}},
{{13'sd4041, 11'sd-874, 13'sd2439}, {12'sd1315, 13'sd-2123, 12'sd1875}, {12'sd1244, 13'sd3039, 13'sd3244}},
{{12'sd-1302, 13'sd-2289, 11'sd-925}, {12'sd1214, 11'sd753, 12'sd-1634}, {10'sd-288, 14'sd-4667, 9'sd230}},
{{9'sd150, 12'sd-1604, 11'sd894}, {12'sd1068, 13'sd3027, 12'sd-1546}, {11'sd-645, 12'sd1238, 13'sd2810}},
{{13'sd2762, 11'sd-656, 13'sd-2215}, {12'sd-1283, 9'sd212, 13'sd-2856}, {11'sd775, 11'sd757, 11'sd830}},
{{11'sd-803, 12'sd1132, 10'sd-383}, {13'sd-2656, 13'sd-2388, 13'sd-2238}, {12'sd1491, 12'sd1689, 9'sd169}},
{{12'sd-1892, 12'sd-1541, 10'sd-296}, {11'sd674, 12'sd-1733, 13'sd2247}, {10'sd-298, 12'sd1139, 13'sd2421}},
{{12'sd1280, 8'sd69, 13'sd-3442}, {12'sd-1158, 12'sd-1631, 9'sd253}, {12'sd1672, 13'sd2057, 13'sd2086}},
{{11'sd-630, 13'sd2143, 10'sd502}, {10'sd443, 12'sd-1918, 13'sd-2231}, {12'sd1638, 10'sd-464, 13'sd-2331}},
{{11'sd641, 12'sd1414, 11'sd-831}, {10'sd346, 13'sd-2120, 13'sd2515}, {13'sd-2130, 13'sd-3648, 8'sd105}},
{{13'sd-3331, 13'sd-3049, 13'sd-2823}, {11'sd898, 10'sd434, 10'sd297}, {13'sd2068, 11'sd568, 11'sd983}},
{{9'sd160, 10'sd409, 7'sd-48}, {12'sd-1373, 12'sd-1609, 12'sd1070}, {13'sd-3169, 13'sd-2235, 12'sd-1227}},
{{9'sd-173, 13'sd-2627, 10'sd-278}, {10'sd415, 13'sd-2639, 9'sd236}, {13'sd3053, 12'sd-1063, 11'sd653}},
{{14'sd-4597, 12'sd-1210, 10'sd317}, {13'sd-2188, 13'sd-2730, 8'sd-67}, {11'sd-956, 10'sd-472, 12'sd1521}},
{{12'sd1174, 9'sd-208, 12'sd-1320}, {8'sd-109, 13'sd2216, 11'sd-831}, {13'sd-2609, 12'sd1342, 7'sd-51}},
{{13'sd-2114, 13'sd2538, 12'sd1072}, {12'sd2047, 13'sd2069, 9'sd143}, {12'sd-1412, 12'sd1551, 12'sd-1417}},
{{14'sd-4324, 13'sd-3467, 9'sd159}, {9'sd-204, 13'sd2273, 8'sd85}, {14'sd-4141, 11'sd-810, 11'sd762}},
{{13'sd4030, 13'sd-2441, 11'sd940}, {14'sd4673, 11'sd837, 13'sd2066}, {12'sd1553, 11'sd734, 12'sd1459}},
{{13'sd3704, 11'sd-757, 13'sd2902}, {12'sd-1153, 11'sd559, 10'sd419}, {12'sd1423, 13'sd2483, 12'sd1454}},
{{11'sd744, 10'sd472, 11'sd-819}, {12'sd-1609, 13'sd2216, 13'sd3099}, {14'sd-4296, 11'sd592, 13'sd3905}},
{{11'sd-983, 12'sd-1299, 13'sd-3882}, {11'sd728, 9'sd-131, 11'sd-524}, {13'sd-2923, 13'sd2049, 12'sd1645}},
{{11'sd-636, 10'sd-271, 9'sd156}, {12'sd-1182, 12'sd1823, 11'sd-514}, {13'sd2242, 9'sd243, 12'sd-1636}},
{{12'sd1029, 13'sd-2170, 11'sd833}, {12'sd1823, 13'sd-2101, 11'sd-972}, {8'sd-86, 11'sd597, 13'sd-2213}},
{{13'sd-3212, 12'sd-1079, 13'sd-2186}, {13'sd2179, 12'sd-1054, 12'sd1161}, {8'sd-83, 12'sd-1603, 11'sd733}},
{{12'sd-1190, 10'sd509, 11'sd594}, {11'sd-526, 12'sd1657, 12'sd-1107}, {12'sd-1343, 12'sd1356, 9'sd-166}},
{{13'sd2815, 12'sd1653, 12'sd-1881}, {11'sd-693, 12'sd1958, 11'sd-671}, {13'sd-2592, 12'sd1429, 12'sd-1693}},
{{5'sd-14, 13'sd2481, 11'sd590}, {12'sd1719, 10'sd-418, 12'sd-1497}, {12'sd-1607, 10'sd303, 8'sd82}},
{{12'sd1882, 12'sd1536, 13'sd3340}, {10'sd-429, 10'sd-492, 13'sd-2865}, {12'sd1887, 13'sd3126, 12'sd1501}},
{{12'sd-1466, 8'sd75, 12'sd-1687}, {13'sd-2054, 11'sd753, 10'sd482}, {13'sd2898, 13'sd-2120, 13'sd-3407}},
{{12'sd-1218, 13'sd-2917, 9'sd-134}, {12'sd-1371, 12'sd1099, 12'sd-1299}, {11'sd-593, 11'sd774, 12'sd1877}},
{{13'sd2992, 10'sd426, 11'sd-902}, {12'sd-1114, 11'sd662, 10'sd346}, {12'sd-1141, 12'sd1817, 12'sd1639}},
{{11'sd-524, 13'sd-2500, 9'sd-202}, {10'sd-509, 13'sd-2375, 10'sd-263}, {12'sd1762, 11'sd-980, 11'sd988}},
{{13'sd-3027, 10'sd427, 12'sd-1769}, {12'sd1611, 12'sd-1673, 12'sd-1549}, {12'sd-1773, 13'sd-2130, 13'sd-3963}}},
{
{{11'sd819, 13'sd2726, 13'sd2860}, {11'sd944, 12'sd-1685, 10'sd490}, {12'sd1043, 13'sd-2203, 13'sd2651}},
{{12'sd1610, 11'sd984, 9'sd226}, {13'sd-3320, 9'sd-245, 13'sd-2357}, {12'sd1137, 12'sd-1257, 9'sd130}},
{{12'sd1224, 10'sd-279, 13'sd-3749}, {8'sd-118, 12'sd-1312, 12'sd-1759}, {13'sd3866, 13'sd2372, 13'sd2289}},
{{13'sd2407, 11'sd-629, 12'sd1288}, {12'sd2017, 12'sd-1189, 13'sd3016}, {10'sd464, 11'sd631, 10'sd261}},
{{13'sd-2329, 13'sd-2342, 12'sd-1934}, {12'sd1759, 13'sd-2426, 10'sd452}, {12'sd-1288, 12'sd1065, 11'sd-821}},
{{13'sd2347, 12'sd1290, 13'sd2664}, {12'sd1030, 12'sd1510, 10'sd491}, {13'sd-3113, 12'sd1448, 13'sd-2393}},
{{13'sd-3858, 10'sd-345, 13'sd-2058}, {10'sd-406, 9'sd234, 13'sd-3738}, {9'sd-208, 14'sd4822, 11'sd-984}},
{{12'sd1258, 11'sd-547, 7'sd59}, {14'sd4174, 13'sd-2290, 13'sd-2156}, {12'sd1538, 12'sd-1690, 12'sd1033}},
{{12'sd-1338, 10'sd-316, 11'sd944}, {10'sd-364, 12'sd1106, 13'sd2579}, {12'sd-1428, 11'sd-768, 12'sd1892}},
{{9'sd225, 11'sd-1023, 13'sd-2910}, {13'sd-2867, 12'sd1810, 12'sd1898}, {12'sd1887, 11'sd580, 12'sd-1942}},
{{8'sd-87, 9'sd251, 12'sd-1418}, {11'sd624, 12'sd-1867, 10'sd-464}, {12'sd-1187, 12'sd-1318, 12'sd1549}},
{{12'sd-1963, 13'sd2750, 13'sd-2169}, {11'sd-719, 11'sd595, 13'sd-2930}, {10'sd434, 13'sd2990, 12'sd-1598}},
{{13'sd-3813, 13'sd-2182, 12'sd-1738}, {13'sd-2449, 12'sd1296, 6'sd25}, {13'sd2201, 12'sd1600, 13'sd2594}},
{{13'sd-3796, 12'sd1432, 11'sd1018}, {12'sd-1080, 11'sd799, 11'sd689}, {12'sd-1139, 12'sd1050, 13'sd-2287}},
{{9'sd236, 12'sd1893, 12'sd-1443}, {11'sd-615, 11'sd652, 13'sd2465}, {13'sd-2383, 12'sd-1757, 11'sd641}},
{{13'sd2360, 11'sd-1001, 11'sd-889}, {12'sd-1047, 12'sd-1893, 13'sd3326}, {13'sd-3229, 11'sd614, 9'sd-180}},
{{12'sd1481, 13'sd2365, 12'sd1916}, {13'sd-2585, 10'sd475, 13'sd-2455}, {13'sd-2722, 11'sd-677, 11'sd-829}},
{{12'sd1994, 12'sd1725, 11'sd797}, {13'sd2290, 13'sd2775, 12'sd1304}, {13'sd-3023, 12'sd1609, 13'sd2658}},
{{13'sd-2499, 12'sd-1073, 13'sd-2414}, {10'sd378, 11'sd-654, 12'sd2013}, {12'sd1589, 12'sd1761, 10'sd370}},
{{13'sd-2504, 12'sd-1509, 12'sd1231}, {12'sd1466, 10'sd341, 13'sd-2364}, {12'sd-1818, 11'sd818, 12'sd-1298}},
{{13'sd-2745, 13'sd-3184, 10'sd-490}, {7'sd-33, 13'sd-2869, 12'sd1256}, {12'sd-1701, 13'sd-2794, 13'sd-3042}},
{{13'sd2773, 12'sd-1157, 10'sd-448}, {11'sd856, 10'sd429, 10'sd-421}, {11'sd589, 9'sd-194, 11'sd549}},
{{12'sd-1798, 11'sd-726, 12'sd1366}, {12'sd-1307, 11'sd689, 12'sd1266}, {12'sd-1812, 13'sd-3354, 11'sd721}},
{{12'sd1847, 12'sd-1755, 12'sd-1515}, {12'sd1377, 12'sd-1971, 13'sd-2298}, {13'sd-2070, 10'sd-326, 12'sd1414}},
{{12'sd-1922, 11'sd-601, 12'sd1499}, {9'sd-160, 13'sd2126, 12'sd-1945}, {13'sd2400, 11'sd-802, 11'sd643}},
{{12'sd-1594, 12'sd1639, 12'sd-1033}, {13'sd2242, 13'sd2205, 11'sd610}, {11'sd536, 11'sd-786, 12'sd1209}},
{{11'sd860, 13'sd-2214, 10'sd-275}, {13'sd2107, 10'sd358, 12'sd1285}, {12'sd-1300, 8'sd70, 12'sd1069}},
{{14'sd-4186, 12'sd1257, 11'sd-633}, {12'sd-1679, 10'sd451, 9'sd-168}, {12'sd1667, 12'sd1770, 13'sd3499}},
{{13'sd-2300, 8'sd-120, 12'sd1445}, {12'sd1173, 13'sd2073, 10'sd-496}, {11'sd1013, 12'sd-1960, 12'sd1899}},
{{13'sd-2389, 13'sd2447, 13'sd2770}, {12'sd1764, 11'sd538, 11'sd-630}, {12'sd-1588, 10'sd-499, 12'sd-1703}},
{{13'sd2614, 12'sd-1791, 13'sd-2161}, {13'sd2143, 13'sd2463, 11'sd528}, {14'sd4913, 14'sd4417, 13'sd2269}},
{{12'sd1698, 13'sd2326, 10'sd-265}, {12'sd2022, 12'sd-1706, 12'sd-1246}, {13'sd2295, 10'sd-303, 12'sd-1812}},
{{13'sd-3729, 13'sd-2509, 12'sd1666}, {12'sd-1967, 12'sd1123, 12'sd1261}, {13'sd4009, 12'sd1098, 11'sd-848}},
{{13'sd-2068, 9'sd-147, 12'sd-1666}, {14'sd-4640, 11'sd744, 12'sd-1694}, {13'sd-3675, 13'sd2112, 11'sd-625}},
{{13'sd2271, 12'sd-1985, 12'sd1823}, {8'sd-80, 12'sd1262, 12'sd-1664}, {13'sd2500, 12'sd-1242, 12'sd-2012}},
{{13'sd-2133, 13'sd2456, 11'sd812}, {12'sd1654, 13'sd-2274, 10'sd-492}, {12'sd1146, 11'sd-515, 12'sd-1973}},
{{13'sd-3019, 10'sd-508, 9'sd-169}, {11'sd908, 12'sd1035, 13'sd-2768}, {11'sd729, 13'sd2473, 9'sd251}},
{{13'sd2870, 11'sd-742, 13'sd-2220}, {12'sd-1050, 12'sd-1481, 12'sd-1558}, {11'sd-826, 12'sd1451, 9'sd-198}},
{{12'sd-1909, 11'sd1013, 11'sd-842}, {13'sd-2334, 12'sd1771, 12'sd-1595}, {12'sd-1990, 10'sd-447, 11'sd936}},
{{11'sd655, 10'sd427, 10'sd-495}, {13'sd2369, 12'sd-1486, 12'sd-2042}, {12'sd-1908, 7'sd48, 11'sd-860}},
{{11'sd-761, 12'sd1418, 12'sd-1365}, {11'sd-769, 11'sd-727, 11'sd829}, {14'sd5108, 11'sd-872, 13'sd2815}},
{{11'sd-763, 8'sd-83, 10'sd490}, {11'sd-987, 12'sd1453, 7'sd44}, {12'sd1348, 13'sd-2474, 12'sd-1931}},
{{12'sd-1746, 13'sd-2244, 12'sd-1643}, {12'sd1273, 12'sd1706, 12'sd-1044}, {12'sd-1857, 11'sd-721, 13'sd2511}},
{{10'sd308, 9'sd213, 11'sd-715}, {9'sd-252, 12'sd2006, 13'sd2297}, {12'sd1853, 10'sd352, 12'sd-1745}},
{{14'sd-4312, 13'sd-3210, 10'sd-460}, {13'sd-2437, 11'sd873, 13'sd-2144}, {13'sd3570, 13'sd3081, 13'sd4002}},
{{13'sd2477, 12'sd-1605, 11'sd-683}, {13'sd2646, 11'sd-726, 12'sd1265}, {13'sd2760, 11'sd-755, 12'sd-1788}},
{{13'sd-2224, 10'sd-420, 12'sd-1773}, {12'sd-1634, 12'sd-1153, 13'sd2714}, {11'sd-538, 11'sd594, 12'sd1888}},
{{8'sd-116, 11'sd-841, 9'sd-154}, {13'sd-4002, 9'sd173, 13'sd-3808}, {12'sd-1374, 11'sd791, 13'sd-2258}},
{{13'sd2613, 13'sd-2482, 12'sd1903}, {4'sd-7, 12'sd-1053, 13'sd-2823}, {13'sd-4053, 11'sd555, 11'sd-541}},
{{11'sd571, 12'sd1142, 13'sd2953}, {7'sd47, 13'sd-2459, 13'sd3295}, {12'sd-1679, 10'sd-272, 13'sd3190}},
{{11'sd569, 13'sd-2366, 12'sd-1314}, {11'sd905, 13'sd-2348, 12'sd1463}, {13'sd2746, 12'sd-1657, 11'sd751}},
{{9'sd-144, 11'sd767, 13'sd-2771}, {10'sd-295, 12'sd-1292, 12'sd-1534}, {12'sd-1231, 9'sd-189, 11'sd618}},
{{11'sd-722, 12'sd1190, 12'sd-1134}, {13'sd2154, 11'sd657, 5'sd-14}, {11'sd-514, 13'sd2275, 11'sd-881}},
{{12'sd1698, 13'sd-3619, 11'sd759}, {13'sd-2064, 10'sd448, 12'sd1493}, {12'sd1960, 11'sd777, 12'sd1912}},
{{10'sd-417, 12'sd-1342, 13'sd-2093}, {12'sd-1699, 12'sd-1046, 13'sd2551}, {12'sd1165, 13'sd2507, 13'sd2958}},
{{12'sd-1672, 12'sd1866, 12'sd-1958}, {13'sd-2333, 11'sd-611, 13'sd2806}, {12'sd-1475, 12'sd1459, 11'sd-946}},
{{12'sd-1654, 12'sd1137, 12'sd-1582}, {10'sd-451, 7'sd-53, 13'sd2136}, {12'sd1263, 11'sd-650, 13'sd-2082}},
{{12'sd-1788, 11'sd594, 12'sd1397}, {13'sd-3433, 11'sd537, 11'sd697}, {8'sd65, 11'sd654, 13'sd3111}},
{{12'sd-1131, 13'sd-2209, 12'sd-1969}, {11'sd-989, 13'sd2711, 13'sd-3017}, {11'sd731, 12'sd-1774, 12'sd1272}},
{{13'sd-2481, 12'sd1283, 13'sd-2829}, {13'sd-3016, 9'sd142, 12'sd-1932}, {13'sd-3789, 12'sd1877, 8'sd-118}},
{{10'sd-464, 12'sd-1674, 13'sd2589}, {12'sd-1626, 12'sd-1150, 13'sd-2895}, {12'sd1139, 12'sd-1030, 7'sd-42}},
{{13'sd2677, 12'sd-1941, 12'sd-1686}, {13'sd2893, 9'sd-180, 12'sd1433}, {11'sd882, 13'sd3748, 11'sd874}},
{{9'sd-246, 13'sd-2187, 13'sd-3189}, {11'sd-573, 11'sd-560, 12'sd1613}, {10'sd-394, 13'sd-2061, 13'sd-2077}},
{{12'sd1403, 12'sd1442, 13'sd2666}, {10'sd387, 13'sd3043, 11'sd899}, {11'sd968, 12'sd-1098, 10'sd275}}},
{
{{11'sd876, 11'sd815, 12'sd1610}, {11'sd-805, 13'sd-2056, 9'sd-167}, {13'sd-2623, 9'sd128, 12'sd-1928}},
{{12'sd1987, 12'sd-1556, 13'sd2134}, {12'sd-2008, 8'sd73, 12'sd-1501}, {13'sd-2855, 10'sd-487, 11'sd743}},
{{14'sd-4503, 10'sd-275, 11'sd-833}, {13'sd-3543, 13'sd2705, 12'sd-1164}, {11'sd873, 8'sd-120, 9'sd132}},
{{11'sd-779, 12'sd-1479, 13'sd-3527}, {12'sd1727, 13'sd3270, 13'sd-2643}, {13'sd2609, 12'sd1903, 12'sd1864}},
{{10'sd425, 13'sd-3052, 13'sd2290}, {8'sd93, 10'sd396, 12'sd1134}, {9'sd192, 9'sd-241, 12'sd-1988}},
{{7'sd-56, 12'sd-1077, 13'sd2326}, {13'sd2208, 12'sd-1436, 12'sd-1820}, {13'sd2256, 13'sd2479, 11'sd626}},
{{13'sd2205, 13'sd2186, 11'sd-901}, {12'sd-1663, 12'sd-1292, 12'sd-1203}, {10'sd474, 8'sd106, 12'sd-1932}},
{{11'sd-935, 13'sd-3525, 13'sd-3010}, {11'sd-783, 12'sd1461, 10'sd455}, {11'sd512, 12'sd1581, 12'sd-1139}},
{{11'sd1022, 13'sd-2335, 12'sd-1144}, {12'sd-1458, 12'sd1468, 12'sd1715}, {13'sd4000, 7'sd55, 10'sd-473}},
{{9'sd-242, 11'sd-977, 10'sd-297}, {12'sd-1189, 13'sd2519, 11'sd755}, {9'sd245, 13'sd-2743, 11'sd-828}},
{{10'sd-411, 12'sd1075, 11'sd706}, {12'sd-1172, 12'sd-1704, 11'sd908}, {12'sd1883, 12'sd-2041, 11'sd-554}},
{{11'sd726, 11'sd872, 13'sd-2293}, {12'sd-1288, 12'sd-1794, 10'sd-454}, {11'sd-1006, 11'sd549, 13'sd-2232}},
{{10'sd-289, 13'sd3024, 13'sd3018}, {12'sd1555, 11'sd614, 11'sd-527}, {12'sd-1504, 13'sd2304, 9'sd-205}},
{{9'sd200, 12'sd-1343, 11'sd843}, {13'sd2381, 12'sd1683, 10'sd429}, {12'sd-1192, 11'sd-1014, 12'sd1571}},
{{11'sd-858, 12'sd-1683, 13'sd-2191}, {13'sd2883, 13'sd2901, 9'sd225}, {12'sd-1126, 12'sd-1268, 9'sd132}},
{{12'sd-1765, 12'sd-1207, 11'sd-884}, {6'sd-31, 12'sd1260, 12'sd1591}, {13'sd2378, 9'sd-231, 13'sd2681}},
{{11'sd903, 12'sd-1049, 11'sd803}, {12'sd1539, 12'sd1187, 13'sd-2491}, {12'sd-1963, 12'sd1440, 12'sd-1260}},
{{14'sd4306, 12'sd-1781, 12'sd-1522}, {13'sd2078, 12'sd-1461, 11'sd670}, {14'sd4536, 8'sd116, 12'sd1306}},
{{11'sd-731, 11'sd-569, 8'sd-110}, {12'sd-1332, 10'sd-479, 12'sd1092}, {10'sd468, 12'sd1076, 12'sd1533}},
{{10'sd-414, 12'sd-1565, 12'sd1791}, {13'sd-2117, 11'sd525, 11'sd751}, {12'sd1456, 13'sd-2443, 12'sd-1782}},
{{13'sd-2742, 12'sd-1301, 12'sd1528}, {11'sd-832, 13'sd2160, 10'sd341}, {12'sd1109, 11'sd548, 11'sd602}},
{{13'sd2214, 11'sd-762, 13'sd-2177}, {13'sd3427, 12'sd-1419, 12'sd-1440}, {12'sd1547, 12'sd1874, 12'sd1574}},
{{11'sd-987, 13'sd2389, 10'sd-343}, {13'sd2507, 12'sd1362, 8'sd81}, {13'sd2088, 11'sd870, 9'sd197}},
{{7'sd-32, 10'sd-465, 12'sd1127}, {11'sd738, 12'sd1937, 6'sd29}, {12'sd-1593, 13'sd2080, 12'sd1782}},
{{12'sd1457, 13'sd2320, 10'sd-298}, {12'sd-1181, 12'sd-1801, 13'sd2081}, {12'sd-1532, 12'sd1768, 12'sd1068}},
{{13'sd2220, 7'sd39, 13'sd2510}, {9'sd144, 10'sd415, 12'sd-1645}, {10'sd373, 11'sd621, 11'sd878}},
{{10'sd-434, 10'sd-313, 11'sd-713}, {12'sd1762, 12'sd-1398, 12'sd-1668}, {11'sd889, 11'sd-921, 10'sd435}},
{{8'sd106, 11'sd1001, 13'sd4043}, {12'sd1141, 11'sd-971, 12'sd-1669}, {12'sd-1062, 12'sd1639, 13'sd2411}},
{{13'sd2189, 12'sd-1076, 13'sd2197}, {8'sd-74, 12'sd1727, 13'sd-2367}, {12'sd1717, 12'sd-1793, 13'sd-2636}},
{{12'sd1667, 12'sd-2018, 12'sd-1587}, {12'sd-1595, 11'sd-695, 10'sd323}, {11'sd845, 13'sd2231, 13'sd2741}},
{{14'sd5966, 11'sd670, 12'sd1177}, {12'sd1247, 11'sd-911, 12'sd-1178}, {8'sd-93, 13'sd-3946, 13'sd-2248}},
{{11'sd-823, 11'sd-572, 12'sd1876}, {13'sd2377, 13'sd-2509, 9'sd219}, {10'sd511, 12'sd1330, 11'sd662}},
{{11'sd578, 11'sd1010, 13'sd2473}, {11'sd596, 12'sd1125, 13'sd2827}, {11'sd687, 13'sd2173, 2'sd1}},
{{12'sd-1302, 13'sd-3581, 13'sd-2991}, {12'sd1619, 12'sd-1235, 10'sd370}, {13'sd2272, 13'sd-2864, 12'sd-1744}},
{{11'sd817, 9'sd-151, 12'sd1988}, {12'sd1333, 13'sd-2843, 12'sd1968}, {11'sd967, 13'sd-2125, 12'sd-1442}},
{{12'sd1342, 13'sd2576, 12'sd-1423}, {11'sd714, 13'sd-2236, 12'sd1664}, {13'sd2265, 13'sd2733, 13'sd2145}},
{{12'sd1238, 12'sd-1192, 13'sd2787}, {12'sd-1398, 12'sd1659, 13'sd2143}, {13'sd-2141, 13'sd-2704, 13'sd-2427}},
{{10'sd481, 12'sd-1580, 13'sd2335}, {12'sd-1177, 11'sd-513, 12'sd1191}, {6'sd23, 13'sd-2288, 12'sd-1101}},
{{11'sd-796, 12'sd-1924, 13'sd-2997}, {9'sd-253, 12'sd1127, 13'sd-2941}, {12'sd1458, 12'sd-1228, 13'sd2659}},
{{13'sd-2543, 13'sd-2110, 13'sd-2660}, {12'sd1414, 12'sd-1066, 11'sd-900}, {13'sd-2571, 12'sd-1465, 12'sd2024}},
{{12'sd1739, 13'sd3194, 13'sd2182}, {12'sd-1552, 11'sd621, 13'sd2493}, {10'sd-366, 11'sd653, 12'sd-1459}},
{{13'sd-3144, 12'sd1614, 12'sd-1552}, {10'sd269, 12'sd1172, 13'sd2607}, {13'sd2226, 13'sd2057, 10'sd473}},
{{9'sd-203, 11'sd517, 12'sd-1135}, {12'sd-1528, 13'sd2675, 12'sd-1884}, {12'sd-1628, 13'sd2247, 8'sd116}},
{{10'sd-289, 12'sd-1629, 13'sd-2335}, {13'sd-2420, 12'sd-1468, 13'sd-2776}, {11'sd941, 9'sd149, 13'sd-2481}},
{{13'sd-2994, 12'sd1786, 10'sd-333}, {13'sd-3324, 10'sd263, 12'sd-1064}, {12'sd-1933, 11'sd-777, 12'sd-1894}},
{{10'sd-328, 13'sd2566, 12'sd-1548}, {6'sd28, 11'sd-935, 12'sd-1162}, {13'sd-2418, 9'sd-220, 12'sd-1907}},
{{12'sd1345, 12'sd1402, 11'sd-531}, {12'sd1556, 11'sd-676, 11'sd584}, {13'sd-2330, 12'sd1993, 12'sd1553}},
{{13'sd-3275, 8'sd-68, 13'sd2291}, {12'sd1380, 12'sd-1660, 13'sd2354}, {13'sd-3306, 11'sd-665, 13'sd2714}},
{{13'sd3647, 12'sd-1685, 13'sd-2168}, {11'sd658, 12'sd1664, 12'sd1309}, {12'sd1622, 13'sd2781, 11'sd-863}},
{{13'sd2425, 12'sd-1567, 11'sd-984}, {11'sd991, 12'sd1120, 13'sd3010}, {11'sd1007, 10'sd469, 13'sd3854}},
{{11'sd-648, 12'sd-1933, 11'sd-664}, {11'sd784, 9'sd-148, 13'sd2917}, {13'sd-2797, 13'sd-2306, 11'sd-642}},
{{12'sd-1499, 9'sd192, 11'sd963}, {11'sd606, 11'sd-737, 12'sd-1173}, {12'sd-1109, 13'sd-2629, 10'sd425}},
{{13'sd-2290, 12'sd1613, 11'sd-1003}, {13'sd2370, 11'sd-650, 12'sd-1728}, {12'sd-1336, 10'sd303, 11'sd685}},
{{13'sd2163, 11'sd732, 12'sd1673}, {13'sd2347, 12'sd1314, 12'sd-1956}, {12'sd1922, 13'sd-2773, 12'sd1531}},
{{12'sd-1257, 12'sd-1902, 13'sd-2358}, {13'sd-2060, 11'sd920, 13'sd-3700}, {12'sd-1341, 10'sd-488, 13'sd-2083}},
{{12'sd-1733, 10'sd-301, 10'sd387}, {13'sd-2120, 12'sd1360, 12'sd1730}, {12'sd-1150, 12'sd1625, 13'sd2422}},
{{11'sd1021, 11'sd852, 11'sd646}, {12'sd-1814, 11'sd-678, 11'sd784}, {12'sd-1742, 13'sd2163, 12'sd-1144}},
{{13'sd-3470, 11'sd869, 11'sd757}, {12'sd-1497, 11'sd977, 12'sd1556}, {12'sd-1965, 11'sd-517, 13'sd3585}},
{{13'sd2231, 12'sd-1213, 13'sd2566}, {9'sd-155, 13'sd2191, 13'sd-2321}, {13'sd-2085, 11'sd-609, 3'sd-3}},
{{12'sd-1747, 11'sd-881, 12'sd-1854}, {13'sd-2988, 13'sd-2591, 13'sd2377}, {13'sd-2134, 13'sd3163, 12'sd1714}},
{{13'sd2749, 12'sd-1062, 12'sd1339}, {12'sd1506, 13'sd-2312, 11'sd-875}, {13'sd2879, 11'sd-675, 13'sd2122}},
{{13'sd2829, 12'sd1836, 11'sd-540}, {13'sd2866, 13'sd-2084, 13'sd-2083}, {7'sd53, 12'sd1696, 11'sd797}},
{{11'sd738, 12'sd-1445, 11'sd683}, {9'sd228, 13'sd2389, 13'sd-2559}, {5'sd-13, 11'sd569, 9'sd147}},
{{13'sd-3245, 12'sd-1438, 13'sd-2245}, {11'sd-530, 11'sd-790, 12'sd1892}, {13'sd-2378, 12'sd-1735, 12'sd1750}}},
{
{{12'sd1395, 13'sd-2803, 12'sd1673}, {12'sd-1535, 12'sd-1913, 10'sd336}, {13'sd-2524, 12'sd-1679, 12'sd2006}},
{{12'sd-1618, 13'sd2138, 12'sd-1541}, {12'sd-1431, 10'sd-405, 13'sd-2244}, {12'sd-1466, 9'sd-156, 13'sd-2123}},
{{10'sd268, 10'sd-336, 11'sd-851}, {12'sd1412, 9'sd-250, 12'sd-1238}, {13'sd2900, 12'sd-1927, 13'sd3342}},
{{11'sd610, 12'sd-1214, 12'sd1308}, {13'sd2234, 11'sd-981, 11'sd987}, {12'sd2006, 11'sd582, 11'sd-827}},
{{11'sd-646, 5'sd-14, 10'sd349}, {12'sd1066, 12'sd-1788, 12'sd1634}, {13'sd2200, 11'sd-523, 10'sd394}},
{{11'sd987, 9'sd160, 12'sd2020}, {11'sd-728, 12'sd-1425, 11'sd-617}, {10'sd288, 13'sd-2433, 12'sd-1394}},
{{12'sd1517, 11'sd519, 12'sd-1431}, {11'sd685, 12'sd-1906, 13'sd-2228}, {11'sd-692, 11'sd996, 12'sd-1026}},
{{11'sd833, 11'sd-965, 12'sd1214}, {13'sd-2157, 13'sd2048, 13'sd2359}, {11'sd-561, 13'sd-2481, 13'sd2103}},
{{12'sd-1837, 7'sd-39, 13'sd-2651}, {12'sd1719, 7'sd37, 11'sd588}, {12'sd1559, 12'sd1501, 10'sd326}},
{{13'sd-2558, 11'sd-934, 12'sd1648}, {8'sd-80, 12'sd-1479, 11'sd-720}, {11'sd-878, 13'sd-2600, 13'sd-2233}},
{{13'sd2321, 11'sd-887, 12'sd1120}, {9'sd173, 13'sd3285, 12'sd-2033}, {11'sd-520, 13'sd2541, 12'sd-1187}},
{{12'sd1497, 12'sd1675, 12'sd2013}, {13'sd-2325, 13'sd-2172, 13'sd-2715}, {12'sd1297, 13'sd-3152, 12'sd-1076}},
{{12'sd-1483, 12'sd-1278, 11'sd-790}, {12'sd-1606, 11'sd-677, 13'sd-2148}, {14'sd-4420, 13'sd-3768, 12'sd-1685}},
{{11'sd-592, 13'sd-2684, 11'sd-660}, {7'sd-41, 13'sd-2495, 11'sd-529}, {13'sd-2578, 12'sd-1880, 13'sd-3057}},
{{13'sd2965, 12'sd1968, 11'sd-517}, {10'sd302, 11'sd-858, 13'sd-2716}, {11'sd-979, 10'sd-462, 13'sd2616}},
{{13'sd2161, 11'sd-880, 13'sd2555}, {12'sd-1483, 10'sd-278, 11'sd-621}, {12'sd1795, 12'sd1469, 13'sd3255}},
{{10'sd472, 11'sd-555, 13'sd-2847}, {12'sd-1725, 13'sd-2843, 12'sd1613}, {11'sd-760, 13'sd2323, 10'sd419}},
{{12'sd-1864, 11'sd-653, 7'sd-40}, {12'sd1122, 13'sd2204, 13'sd3395}, {13'sd-2114, 13'sd3660, 13'sd2497}},
{{11'sd1000, 12'sd1554, 10'sd-316}, {13'sd-2316, 13'sd-3022, 12'sd-1490}, {12'sd-1798, 12'sd1457, 13'sd2062}},
{{10'sd-511, 11'sd-733, 11'sd-983}, {11'sd-629, 13'sd3069, 13'sd2935}, {13'sd2096, 12'sd-1121, 12'sd1863}},
{{12'sd1032, 13'sd-2827, 11'sd585}, {12'sd1437, 11'sd-544, 12'sd1618}, {12'sd-1746, 13'sd-2463, 13'sd-2495}},
{{13'sd-2558, 13'sd-3167, 10'sd354}, {9'sd236, 10'sd426, 11'sd803}, {12'sd1265, 12'sd-1999, 10'sd424}},
{{11'sd689, 9'sd236, 12'sd-1123}, {13'sd2353, 10'sd462, 13'sd-2297}, {12'sd1216, 11'sd900, 10'sd394}},
{{6'sd16, 12'sd-2035, 13'sd2184}, {12'sd-1374, 12'sd1388, 12'sd1558}, {12'sd-1301, 10'sd409, 12'sd-1640}},
{{12'sd1206, 13'sd2889, 10'sd296}, {13'sd-2250, 13'sd2631, 12'sd1248}, {10'sd341, 13'sd3025, 13'sd2116}},
{{13'sd2153, 12'sd-1153, 12'sd1412}, {13'sd3015, 12'sd1866, 12'sd-1786}, {13'sd2522, 12'sd1118, 12'sd-1663}},
{{13'sd-2942, 12'sd-1393, 11'sd734}, {12'sd-1933, 11'sd775, 11'sd804}, {12'sd-1723, 12'sd1555, 11'sd609}},
{{11'sd956, 11'sd886, 12'sd-1587}, {10'sd469, 12'sd1125, 12'sd-1699}, {12'sd1789, 11'sd850, 10'sd287}},
{{12'sd1594, 12'sd1958, 11'sd-679}, {12'sd1344, 11'sd-676, 11'sd738}, {12'sd1358, 13'sd-2159, 11'sd1019}},
{{12'sd1942, 12'sd1908, 12'sd-1533}, {12'sd1603, 12'sd-1042, 13'sd-2672}, {12'sd1244, 13'sd2051, 8'sd106}},
{{11'sd984, 7'sd58, 11'sd-748}, {13'sd-2248, 13'sd2859, 11'sd971}, {9'sd176, 13'sd2526, 13'sd2682}},
{{11'sd-768, 11'sd-745, 12'sd1050}, {12'sd-1271, 10'sd-468, 12'sd-1172}, {9'sd-172, 12'sd-1776, 11'sd548}},
{{10'sd508, 12'sd1165, 12'sd-1925}, {13'sd-2269, 9'sd-168, 13'sd2365}, {13'sd-2181, 11'sd-586, 12'sd1406}},
{{9'sd253, 12'sd-1674, 10'sd-277}, {11'sd-813, 11'sd-514, 13'sd2647}, {13'sd3957, 12'sd1791, 13'sd2171}},
{{12'sd1639, 12'sd1404, 11'sd-884}, {11'sd-557, 13'sd2050, 12'sd-1456}, {13'sd-2811, 13'sd-2763, 10'sd477}},
{{11'sd-903, 13'sd-2083, 10'sd-471}, {9'sd-161, 11'sd796, 11'sd-783}, {13'sd2397, 13'sd-2313, 13'sd-2119}},
{{13'sd-2068, 12'sd-1248, 12'sd-1128}, {12'sd-1785, 12'sd-1502, 10'sd353}, {12'sd-1727, 11'sd-831, 13'sd-2316}},
{{12'sd1245, 13'sd2377, 13'sd-2180}, {12'sd-2015, 12'sd1042, 11'sd699}, {13'sd-2641, 11'sd-940, 10'sd-361}},
{{11'sd1013, 12'sd-1669, 10'sd-378}, {12'sd1273, 13'sd2365, 10'sd286}, {11'sd520, 13'sd-2189, 13'sd2792}},
{{12'sd1447, 12'sd-1027, 10'sd435}, {13'sd-2473, 12'sd-1413, 12'sd1649}, {13'sd-2173, 9'sd-247, 11'sd1008}},
{{11'sd577, 10'sd257, 13'sd-2594}, {13'sd-2284, 13'sd-3432, 12'sd-1132}, {10'sd-340, 13'sd-4086, 11'sd737}},
{{10'sd476, 12'sd1491, 10'sd-351}, {12'sd1374, 10'sd-483, 12'sd1629}, {12'sd1080, 12'sd-1766, 12'sd-1420}},
{{10'sd276, 12'sd-1798, 13'sd2401}, {13'sd2717, 12'sd1911, 11'sd-613}, {11'sd-662, 12'sd1782, 12'sd-1608}},
{{8'sd-103, 11'sd1007, 12'sd1724}, {11'sd563, 8'sd93, 12'sd1907}, {9'sd-216, 13'sd2846, 10'sd318}},
{{10'sd340, 8'sd96, 13'sd2079}, {11'sd518, 13'sd-2118, 12'sd1302}, {13'sd2320, 13'sd-2470, 12'sd1456}},
{{12'sd1823, 9'sd-178, 12'sd2041}, {12'sd1787, 13'sd2923, 11'sd562}, {13'sd2485, 10'sd-332, 12'sd1430}},
{{13'sd2528, 13'sd2633, 12'sd1367}, {13'sd-2199, 13'sd-2152, 12'sd-1295}, {13'sd-2057, 13'sd2571, 13'sd2943}},
{{13'sd-2264, 13'sd-3218, 12'sd1136}, {12'sd1271, 5'sd-13, 10'sd396}, {12'sd1326, 12'sd-1684, 7'sd34}},
{{11'sd-716, 13'sd2256, 12'sd-1292}, {12'sd-1761, 11'sd-979, 12'sd-1666}, {11'sd732, 13'sd2111, 12'sd-1673}},
{{13'sd-2839, 12'sd1374, 12'sd-1402}, {9'sd138, 8'sd84, 8'sd106}, {10'sd-475, 13'sd3360, 11'sd600}},
{{12'sd-1807, 12'sd1094, 10'sd-379}, {11'sd-655, 11'sd-981, 11'sd789}, {12'sd1335, 10'sd-416, 12'sd-1953}},
{{12'sd1070, 13'sd2113, 11'sd571}, {13'sd-2085, 12'sd1513, 12'sd1298}, {8'sd87, 11'sd847, 13'sd-2314}},
{{12'sd1598, 13'sd-2301, 11'sd-895}, {12'sd1647, 13'sd2264, 13'sd2274}, {10'sd-369, 13'sd2515, 12'sd-1211}},
{{13'sd2345, 11'sd771, 12'sd1195}, {13'sd-2449, 11'sd-938, 10'sd-429}, {13'sd-2948, 11'sd-976, 12'sd1495}},
{{13'sd-3549, 9'sd220, 6'sd-29}, {13'sd-2853, 11'sd-1021, 13'sd2986}, {11'sd-642, 13'sd-2939, 13'sd-2562}},
{{12'sd-1615, 13'sd2567, 12'sd1903}, {12'sd-2000, 12'sd2036, 13'sd-2068}, {13'sd2444, 13'sd-2274, 11'sd-543}},
{{11'sd874, 13'sd-2615, 10'sd-340}, {13'sd-2940, 12'sd1223, 11'sd-817}, {13'sd-2441, 11'sd977, 11'sd984}},
{{12'sd1506, 13'sd-2056, 13'sd2691}, {12'sd1390, 10'sd256, 8'sd91}, {10'sd-433, 6'sd31, 11'sd883}},
{{11'sd984, 13'sd2190, 12'sd1100}, {10'sd-473, 11'sd985, 13'sd-2561}, {12'sd-1291, 12'sd-1470, 13'sd-2678}},
{{11'sd-975, 13'sd-3049, 11'sd535}, {13'sd2450, 11'sd-790, 12'sd1559}, {12'sd-1425, 12'sd-1588, 10'sd-467}},
{{12'sd-1330, 12'sd-1767, 11'sd-822}, {12'sd1400, 12'sd-1240, 11'sd-875}, {11'sd515, 12'sd1745, 9'sd-228}},
{{13'sd2241, 11'sd732, 9'sd-170}, {12'sd-1144, 13'sd2463, 12'sd1666}, {12'sd1853, 9'sd166, 12'sd1392}},
{{12'sd1223, 10'sd-321, 12'sd-1801}, {11'sd732, 13'sd-2347, 13'sd2848}, {11'sd-713, 11'sd-829, 12'sd-1946}},
{{12'sd1395, 12'sd1283, 12'sd-1309}, {12'sd1116, 13'sd2711, 11'sd911}, {12'sd-1629, 12'sd-1230, 13'sd-2110}}},
{
{{12'sd1676, 2'sd1, 10'sd289}, {11'sd-739, 12'sd-2035, 12'sd1772}, {10'sd258, 13'sd2613, 11'sd-563}},
{{12'sd-1581, 10'sd290, 11'sd512}, {11'sd753, 8'sd81, 10'sd257}, {12'sd-1205, 10'sd-454, 13'sd-3327}},
{{12'sd-1085, 8'sd-109, 10'sd447}, {13'sd3359, 11'sd-949, 12'sd-1401}, {13'sd2125, 13'sd2774, 12'sd-1411}},
{{12'sd-1809, 12'sd2020, 12'sd1139}, {7'sd-56, 12'sd1564, 13'sd-2341}, {13'sd-3254, 12'sd-1463, 13'sd-2683}},
{{10'sd-322, 12'sd-1874, 12'sd-1519}, {13'sd2106, 12'sd1600, 12'sd-1559}, {12'sd-1380, 13'sd-2657, 12'sd-1572}},
{{12'sd-1131, 9'sd-184, 12'sd-1813}, {10'sd407, 12'sd-1888, 12'sd1566}, {12'sd1946, 13'sd-2520, 13'sd-2245}},
{{13'sd-2667, 12'sd-1726, 12'sd1824}, {8'sd99, 11'sd-787, 10'sd297}, {10'sd405, 13'sd2548, 11'sd-681}},
{{11'sd653, 12'sd-1692, 13'sd-2079}, {13'sd3801, 11'sd562, 14'sd-4574}, {13'sd2631, 11'sd-843, 12'sd-1499}},
{{13'sd3687, 14'sd4556, 10'sd-443}, {12'sd-1458, 11'sd-914, 11'sd982}, {11'sd-642, 10'sd353, 13'sd-3088}},
{{12'sd1726, 13'sd2632, 13'sd2653}, {13'sd-2208, 13'sd2627, 13'sd-2302}, {12'sd-1219, 12'sd1315, 13'sd2240}},
{{12'sd-1893, 12'sd1166, 13'sd-2513}, {13'sd2049, 13'sd-2718, 13'sd-2480}, {13'sd-2130, 13'sd-2541, 11'sd585}},
{{10'sd294, 12'sd1416, 12'sd-1627}, {13'sd-2822, 12'sd1595, 12'sd-1053}, {12'sd1787, 12'sd-1367, 12'sd1848}},
{{9'sd225, 12'sd-1545, 12'sd-1725}, {12'sd1573, 12'sd-1136, 12'sd1119}, {14'sd4485, 14'sd5814, 13'sd3003}},
{{9'sd-230, 12'sd-1635, 11'sd931}, {12'sd-1130, 12'sd-1186, 7'sd-52}, {12'sd1770, 12'sd-2021, 13'sd-2865}},
{{6'sd23, 12'sd-1495, 13'sd-2476}, {12'sd-1938, 13'sd2107, 13'sd-2217}, {13'sd-2051, 12'sd-1871, 13'sd-3962}},
{{12'sd-1932, 12'sd-1042, 12'sd-1265}, {12'sd1260, 12'sd1493, 12'sd-1304}, {10'sd329, 13'sd-2262, 10'sd-312}},
{{12'sd-1714, 11'sd520, 12'sd1912}, {13'sd2309, 12'sd-1730, 11'sd947}, {12'sd1337, 12'sd1474, 12'sd1287}},
{{13'sd3363, 11'sd-526, 11'sd884}, {13'sd3813, 12'sd-1128, 12'sd1256}, {13'sd3228, 11'sd-1022, 12'sd1533}},
{{11'sd-518, 11'sd-761, 12'sd-1053}, {12'sd-1321, 13'sd-2393, 12'sd-1892}, {10'sd-379, 11'sd-984, 13'sd-3341}},
{{13'sd2333, 13'sd-2628, 11'sd-771}, {13'sd-2805, 13'sd-2817, 13'sd-2923}, {12'sd2033, 13'sd2213, 10'sd-499}},
{{14'sd4609, 13'sd2111, 12'sd1964}, {11'sd683, 10'sd393, 12'sd1785}, {13'sd2848, 11'sd675, 12'sd-1815}},
{{12'sd1499, 9'sd-168, 13'sd2433}, {11'sd-977, 11'sd846, 10'sd344}, {11'sd-969, 12'sd1285, 10'sd-434}},
{{13'sd3117, 11'sd-853, 13'sd-2836}, {13'sd-2090, 11'sd-828, 13'sd-2683}, {9'sd145, 12'sd-1451, 12'sd-1973}},
{{13'sd-2227, 12'sd-1139, 11'sd743}, {12'sd1635, 11'sd-685, 13'sd-3167}, {9'sd248, 13'sd-2895, 11'sd-752}},
{{11'sd714, 13'sd-2641, 10'sd-357}, {10'sd409, 11'sd-829, 12'sd1809}, {12'sd-1396, 11'sd660, 12'sd1881}},
{{13'sd-3087, 8'sd102, 11'sd909}, {13'sd-2723, 10'sd-440, 11'sd-899}, {13'sd-2366, 13'sd-2638, 12'sd-1602}},
{{13'sd2240, 12'sd-1392, 13'sd-2530}, {10'sd-500, 12'sd1750, 13'sd2267}, {12'sd-1246, 11'sd-873, 12'sd-1046}},
{{12'sd-1629, 11'sd760, 10'sd401}, {12'sd-1160, 12'sd-1448, 13'sd2278}, {13'sd-3036, 11'sd-598, 12'sd-1925}},
{{9'sd179, 11'sd989, 13'sd-2379}, {12'sd1502, 12'sd1208, 10'sd510}, {11'sd649, 10'sd336, 13'sd2398}},
{{12'sd-1972, 10'sd443, 13'sd2183}, {12'sd-1258, 11'sd-575, 13'sd3006}, {12'sd-1993, 13'sd-3088, 11'sd888}},
{{11'sd-873, 10'sd-509, 13'sd-4002}, {13'sd2380, 13'sd-3270, 11'sd538}, {13'sd2486, 12'sd1428, 12'sd-1105}},
{{11'sd710, 10'sd-319, 11'sd1016}, {12'sd1451, 13'sd2587, 12'sd1834}, {13'sd-2774, 11'sd723, 11'sd-834}},
{{13'sd-2447, 11'sd-904, 12'sd-1676}, {11'sd-655, 9'sd194, 9'sd195}, {13'sd-2239, 12'sd1684, 10'sd-498}},
{{10'sd277, 11'sd-678, 13'sd-2363}, {13'sd-3723, 10'sd272, 9'sd212}, {13'sd-3551, 11'sd-694, 13'sd-3006}},
{{12'sd-1255, 13'sd-2224, 13'sd2500}, {8'sd-97, 13'sd-2448, 11'sd873}, {12'sd1916, 12'sd-1171, 10'sd503}},
{{12'sd-1063, 12'sd-2022, 12'sd-1290}, {11'sd-1012, 13'sd-2173, 13'sd-2182}, {12'sd1221, 12'sd2028, 12'sd1911}},
{{12'sd-1233, 13'sd2445, 11'sd853}, {10'sd-413, 13'sd2369, 12'sd-1306}, {12'sd-1119, 11'sd622, 13'sd-2515}},
{{11'sd-661, 13'sd2108, 11'sd-522}, {13'sd-2821, 12'sd1928, 11'sd-520}, {11'sd-816, 10'sd-315, 12'sd-1586}},
{{12'sd1468, 12'sd1392, 13'sd2981}, {13'sd-2359, 11'sd774, 13'sd3159}, {13'sd-2221, 12'sd1773, 13'sd3001}},
{{13'sd-2615, 12'sd1757, 11'sd-949}, {13'sd-3064, 13'sd2302, 12'sd1313}, {14'sd-4152, 13'sd-3136, 12'sd-1134}},
{{13'sd-2933, 10'sd464, 12'sd1882}, {12'sd-1954, 13'sd2840, 12'sd-1544}, {7'sd52, 14'sd4344, 12'sd1091}},
{{13'sd-2196, 13'sd2330, 11'sd-917}, {13'sd-2583, 12'sd1482, 13'sd3363}, {12'sd1451, 14'sd5230, 14'sd5794}},
{{12'sd-1915, 12'sd-1143, 12'sd1240}, {11'sd928, 12'sd1832, 13'sd2189}, {13'sd2755, 10'sd-405, 11'sd876}},
{{13'sd2469, 13'sd2086, 12'sd-1725}, {12'sd1611, 13'sd-2542, 13'sd2202}, {13'sd2519, 9'sd-250, 13'sd2864}},
{{12'sd1947, 13'sd-2548, 12'sd1712}, {10'sd334, 11'sd-964, 13'sd2263}, {13'sd-2297, 9'sd-160, 10'sd-482}},
{{10'sd292, 12'sd-1229, 13'sd2131}, {12'sd1991, 12'sd-1435, 11'sd1004}, {12'sd1318, 12'sd1815, 13'sd2935}},
{{12'sd-1856, 13'sd2841, 12'sd-1658}, {12'sd1777, 10'sd500, 13'sd2321}, {12'sd-1035, 9'sd-210, 13'sd2518}},
{{10'sd473, 5'sd11, 13'sd-2505}, {13'sd-3684, 11'sd-670, 13'sd-2129}, {11'sd760, 14'sd4309, 13'sd2560}},
{{14'sd4538, 13'sd2403, 12'sd1595}, {13'sd2133, 11'sd995, 13'sd-3172}, {13'sd2656, 13'sd-2465, 8'sd-114}},
{{13'sd2087, 12'sd-1234, 11'sd-781}, {11'sd738, 11'sd671, 11'sd908}, {13'sd-3434, 14'sd-4617, 13'sd-3611}},
{{13'sd-3590, 5'sd11, 12'sd1042}, {12'sd-1889, 12'sd-1923, 11'sd-761}, {11'sd-951, 11'sd620, 12'sd-1856}},
{{13'sd-2833, 9'sd174, 12'sd-1046}, {13'sd2094, 11'sd-704, 12'sd-1877}, {10'sd-261, 12'sd1268, 12'sd2029}},
{{13'sd-2222, 11'sd-541, 13'sd2051}, {7'sd-53, 13'sd2072, 13'sd2870}, {13'sd-2268, 12'sd1433, 9'sd-176}},
{{11'sd-816, 12'sd-1457, 12'sd-1380}, {13'sd3051, 12'sd-1531, 13'sd-2797}, {6'sd22, 12'sd-1235, 11'sd758}},
{{13'sd-2252, 13'sd-2227, 10'sd380}, {10'sd428, 13'sd2355, 13'sd2164}, {12'sd1299, 13'sd2115, 12'sd1662}},
{{11'sd-792, 11'sd-647, 12'sd1683}, {11'sd911, 12'sd1526, 11'sd788}, {10'sd-315, 10'sd-451, 12'sd1970}},
{{10'sd478, 11'sd-918, 13'sd-2496}, {10'sd-471, 13'sd-2789, 13'sd-2750}, {13'sd-2300, 13'sd-2405, 11'sd-855}},
{{11'sd-579, 12'sd1574, 13'sd-3250}, {8'sd82, 10'sd317, 12'sd-1090}, {11'sd-784, 13'sd-4052, 14'sd-5581}},
{{13'sd-2543, 12'sd-1373, 12'sd1433}, {13'sd-2566, 10'sd-495, 11'sd-522}, {13'sd2404, 11'sd-921, 9'sd-241}},
{{12'sd-2022, 13'sd2244, 13'sd2219}, {13'sd2438, 13'sd2610, 13'sd2239}, {12'sd1679, 13'sd2552, 14'sd5786}},
{{12'sd-1765, 12'sd-1692, 11'sd881}, {4'sd7, 10'sd-370, 13'sd-2726}, {12'sd-1069, 11'sd527, 10'sd444}},
{{13'sd-2139, 10'sd-494, 13'sd-2822}, {12'sd1370, 9'sd137, 13'sd-3103}, {12'sd-1369, 13'sd-2965, 11'sd-764}},
{{13'sd-2828, 13'sd-3546, 12'sd-1164}, {12'sd-1982, 13'sd-2564, 11'sd-761}, {8'sd-115, 11'sd-531, 13'sd3751}},
{{12'sd-1242, 13'sd2090, 10'sd-411}, {12'sd-1816, 10'sd-500, 11'sd-536}, {10'sd-272, 12'sd-1844, 12'sd1393}}},
{
{{11'sd863, 13'sd-2489, 12'sd1984}, {13'sd-2462, 11'sd-713, 12'sd1734}, {10'sd-504, 13'sd-2682, 10'sd278}},
{{13'sd-2452, 12'sd-1905, 11'sd1012}, {13'sd2373, 13'sd2254, 7'sd-56}, {12'sd-1228, 12'sd-1927, 11'sd-926}},
{{11'sd858, 8'sd-78, 11'sd-603}, {13'sd-2263, 10'sd396, 12'sd-1805}, {14'sd-4943, 13'sd-3923, 12'sd-1778}},
{{9'sd248, 12'sd-1074, 13'sd2063}, {12'sd-1619, 13'sd-2170, 13'sd-2491}, {12'sd1529, 12'sd1299, 12'sd1456}},
{{12'sd2034, 13'sd-2245, 6'sd-22}, {11'sd-578, 12'sd-1347, 12'sd1150}, {11'sd-952, 12'sd1077, 11'sd753}},
{{11'sd-907, 10'sd479, 13'sd-2991}, {12'sd1330, 13'sd-2236, 8'sd-113}, {10'sd319, 13'sd-2579, 10'sd291}},
{{12'sd-1195, 11'sd-886, 10'sd-472}, {11'sd-723, 12'sd1205, 12'sd1212}, {14'sd4262, 13'sd2636, 10'sd-505}},
{{11'sd-894, 12'sd1198, 10'sd499}, {12'sd-1510, 12'sd-1102, 13'sd-3054}, {13'sd-2185, 10'sd-362, 13'sd-3610}},
{{9'sd-159, 12'sd1268, 13'sd-2158}, {13'sd-2155, 11'sd-583, 13'sd-2444}, {11'sd757, 13'sd2108, 13'sd-2107}},
{{13'sd2703, 13'sd2179, 13'sd2431}, {10'sd-366, 10'sd-263, 12'sd1506}, {13'sd2751, 11'sd812, 12'sd1416}},
{{10'sd-394, 12'sd-1134, 13'sd2312}, {10'sd398, 9'sd145, 11'sd-801}, {12'sd1458, 12'sd1129, 11'sd642}},
{{9'sd243, 12'sd-1731, 12'sd1716}, {13'sd-2715, 12'sd1283, 12'sd-1295}, {12'sd1976, 12'sd-1763, 12'sd1603}},
{{10'sd282, 12'sd-1385, 11'sd-612}, {13'sd2623, 7'sd-62, 12'sd-1757}, {12'sd-1266, 8'sd102, 13'sd-3730}},
{{12'sd-1401, 12'sd-1319, 13'sd-2264}, {12'sd-1413, 12'sd-1396, 10'sd329}, {13'sd-2273, 12'sd2041, 7'sd-55}},
{{10'sd510, 10'sd-492, 12'sd-1194}, {13'sd2849, 8'sd-88, 8'sd-67}, {9'sd-239, 12'sd-1267, 13'sd-3691}},
{{10'sd324, 12'sd-1614, 11'sd-615}, {12'sd-1604, 11'sd698, 13'sd-2049}, {11'sd-838, 12'sd1501, 11'sd725}},
{{13'sd2639, 13'sd2383, 12'sd1804}, {13'sd3070, 13'sd2516, 13'sd-2549}, {13'sd3244, 10'sd352, 12'sd-1331}},
{{12'sd1071, 7'sd55, 11'sd769}, {12'sd1543, 13'sd-2809, 10'sd442}, {13'sd-3268, 12'sd1412, 12'sd1150}},
{{12'sd1744, 13'sd2609, 13'sd2411}, {11'sd796, 12'sd1878, 12'sd-1044}, {12'sd1509, 11'sd519, 9'sd244}},
{{12'sd1231, 12'sd-1560, 10'sd350}, {12'sd-1368, 13'sd2441, 11'sd-585}, {11'sd-912, 12'sd-1338, 13'sd2406}},
{{8'sd92, 13'sd-2058, 13'sd2292}, {12'sd1280, 12'sd-1374, 5'sd-14}, {12'sd-1417, 12'sd-1592, 11'sd-670}},
{{11'sd901, 13'sd-3058, 12'sd1153}, {11'sd801, 12'sd-1912, 13'sd-2682}, {9'sd130, 10'sd-455, 13'sd-3071}},
{{12'sd-1921, 13'sd2647, 13'sd-3038}, {11'sd-730, 12'sd-1932, 12'sd-1124}, {10'sd-499, 11'sd570, 12'sd1765}},
{{13'sd2096, 12'sd-1254, 13'sd-3247}, {10'sd344, 12'sd1653, 13'sd-2308}, {13'sd2666, 7'sd-34, 12'sd-1025}},
{{12'sd1412, 12'sd-1378, 12'sd-1044}, {12'sd-1897, 13'sd2566, 12'sd1564}, {11'sd-811, 13'sd-2413, 13'sd2890}},
{{11'sd-816, 13'sd2100, 8'sd-72}, {10'sd434, 13'sd-2459, 11'sd-990}, {12'sd-1154, 11'sd-541, 12'sd1587}},
{{12'sd1613, 11'sd-634, 12'sd-1298}, {13'sd2250, 12'sd1875, 12'sd-1154}, {12'sd1951, 11'sd648, 12'sd-2022}},
{{13'sd2125, 13'sd-2248, 9'sd-165}, {12'sd1530, 11'sd-613, 11'sd-723}, {9'sd-180, 13'sd2733, 13'sd-2194}},
{{11'sd-562, 13'sd-2294, 10'sd-424}, {9'sd-220, 13'sd-2406, 13'sd2215}, {12'sd1901, 8'sd116, 11'sd-670}},
{{12'sd-1638, 6'sd-29, 13'sd-2329}, {10'sd474, 9'sd-140, 13'sd2069}, {13'sd-2355, 11'sd-622, 11'sd622}},
{{13'sd-2318, 12'sd-1733, 13'sd-2058}, {12'sd-1147, 11'sd1009, 13'sd-2647}, {12'sd1535, 10'sd373, 8'sd104}},
{{10'sd286, 13'sd2792, 13'sd-2641}, {10'sd439, 13'sd-2403, 11'sd1002}, {13'sd-2691, 11'sd-949, 13'sd-2872}},
{{8'sd-72, 12'sd1138, 13'sd2780}, {11'sd-686, 13'sd-2155, 9'sd-145}, {10'sd362, 11'sd-911, 12'sd1286}},
{{12'sd-1282, 9'sd139, 11'sd915}, {11'sd-863, 12'sd1403, 12'sd2024}, {13'sd2788, 12'sd1790, 11'sd939}},
{{12'sd1498, 13'sd-2239, 12'sd1898}, {12'sd-1306, 11'sd654, 13'sd3039}, {13'sd2519, 13'sd-2379, 9'sd210}},
{{9'sd213, 9'sd192, 12'sd-1213}, {12'sd1917, 10'sd304, 13'sd2384}, {12'sd1130, 11'sd-573, 13'sd2468}},
{{12'sd1460, 13'sd-2531, 7'sd-61}, {10'sd-273, 13'sd2120, 10'sd-500}, {12'sd1977, 13'sd2664, 10'sd-504}},
{{12'sd1233, 12'sd1039, 13'sd2081}, {12'sd-1200, 12'sd-1425, 13'sd2115}, {12'sd1922, 13'sd-2238, 12'sd1995}},
{{6'sd26, 12'sd-1891, 12'sd1695}, {12'sd-1566, 12'sd1101, 12'sd1176}, {11'sd954, 12'sd-1627, 11'sd-802}},
{{13'sd-2068, 7'sd-34, 11'sd-636}, {8'sd-96, 8'sd-94, 13'sd-2500}, {12'sd1339, 13'sd-2273, 11'sd-531}},
{{12'sd1841, 13'sd-2826, 13'sd-3112}, {12'sd1762, 12'sd-1530, 10'sd499}, {10'sd-466, 11'sd873, 12'sd-1290}},
{{12'sd-1559, 13'sd2813, 12'sd1308}, {6'sd24, 12'sd-1920, 9'sd146}, {12'sd-1645, 13'sd-3504, 12'sd-1167}},
{{11'sd-794, 12'sd1556, 12'sd-1802}, {12'sd1701, 10'sd360, 12'sd1518}, {12'sd1211, 12'sd-1111, 13'sd2084}},
{{11'sd-581, 11'sd-987, 13'sd2785}, {12'sd-1677, 13'sd-2241, 13'sd-2278}, {11'sd731, 13'sd2388, 12'sd-1540}},
{{8'sd-98, 12'sd-1846, 13'sd2214}, {12'sd1833, 12'sd1138, 10'sd434}, {12'sd-1143, 13'sd2051, 11'sd-653}},
{{11'sd-682, 12'sd-1601, 10'sd363}, {10'sd377, 8'sd-97, 12'sd1127}, {12'sd-1751, 12'sd-1537, 13'sd-2579}},
{{10'sd-455, 11'sd864, 12'sd1940}, {12'sd1903, 13'sd-2201, 12'sd-1460}, {11'sd-948, 9'sd242, 11'sd-709}},
{{13'sd2549, 12'sd1193, 13'sd2681}, {9'sd184, 11'sd-769, 13'sd-2419}, {12'sd-1365, 13'sd-3411, 8'sd100}},
{{11'sd1020, 12'sd-1350, 13'sd-2495}, {12'sd-1639, 8'sd-113, 12'sd1367}, {11'sd856, 11'sd754, 12'sd-1622}},
{{13'sd-3035, 9'sd-165, 12'sd-1072}, {11'sd875, 13'sd2494, 10'sd469}, {11'sd-728, 13'sd2351, 11'sd811}},
{{13'sd-2748, 10'sd509, 10'sd425}, {12'sd-1404, 11'sd859, 12'sd1816}, {10'sd341, 12'sd-1769, 11'sd614}},
{{13'sd2896, 10'sd-392, 13'sd-2591}, {10'sd503, 12'sd1246, 13'sd-2466}, {11'sd621, 12'sd-1381, 12'sd1889}},
{{13'sd-2517, 12'sd1951, 8'sd112}, {10'sd475, 5'sd-11, 11'sd1017}, {11'sd952, 8'sd88, 9'sd248}},
{{13'sd-2329, 11'sd541, 11'sd-600}, {10'sd299, 8'sd125, 12'sd-1325}, {12'sd1864, 2'sd-1, 7'sd62}},
{{9'sd-174, 12'sd-1255, 13'sd3606}, {12'sd-1133, 12'sd1461, 13'sd3512}, {13'sd-3371, 13'sd-2621, 13'sd-2463}},
{{11'sd716, 12'sd1904, 12'sd-1420}, {13'sd2123, 13'sd-2349, 9'sd222}, {13'sd-2524, 12'sd-1486, 11'sd773}},
{{10'sd-355, 11'sd568, 11'sd589}, {12'sd-1093, 12'sd-1618, 11'sd-1022}, {13'sd-4029, 13'sd-2299, 10'sd-396}},
{{10'sd454, 11'sd-865, 13'sd-2234}, {13'sd2898, 11'sd-1015, 12'sd1927}, {13'sd2120, 11'sd736, 12'sd-1952}},
{{12'sd-1638, 12'sd-1977, 13'sd2299}, {9'sd-133, 12'sd-1160, 12'sd-1232}, {10'sd-394, 9'sd-246, 13'sd3622}},
{{11'sd-803, 11'sd866, 10'sd-370}, {13'sd2341, 12'sd1375, 10'sd368}, {13'sd2441, 10'sd511, 12'sd1711}},
{{12'sd1449, 12'sd1949, 13'sd-2376}, {12'sd-1169, 9'sd-179, 13'sd-2281}, {12'sd1095, 8'sd65, 13'sd2200}},
{{12'sd-1867, 12'sd1733, 11'sd-972}, {12'sd-1909, 12'sd-1559, 11'sd737}, {9'sd142, 11'sd-756, 10'sd-480}},
{{11'sd-997, 13'sd3259, 13'sd2344}, {13'sd-2996, 12'sd-1654, 11'sd591}, {12'sd-1702, 13'sd2405, 13'sd2718}},
{{12'sd2033, 13'sd-2809, 10'sd-475}, {12'sd1361, 12'sd-1650, 12'sd1312}, {13'sd-2828, 10'sd-369, 13'sd-2390}}},
{
{{12'sd1394, 11'sd-657, 11'sd-938}, {11'sd-941, 12'sd1996, 13'sd-2329}, {13'sd-3505, 13'sd-2444, 12'sd1462}},
{{13'sd2550, 12'sd1738, 12'sd1321}, {10'sd-327, 11'sd-721, 11'sd-536}, {13'sd2615, 12'sd-1064, 12'sd-1555}},
{{12'sd-1777, 13'sd-2790, 13'sd-3109}, {13'sd2418, 12'sd-1537, 11'sd871}, {7'sd-38, 13'sd-3182, 13'sd-2408}},
{{13'sd3634, 13'sd3847, 10'sd435}, {9'sd-180, 12'sd-1099, 13'sd2052}, {10'sd-438, 8'sd-71, 10'sd-361}},
{{10'sd298, 12'sd1226, 12'sd-1033}, {13'sd3320, 12'sd1814, 13'sd-2422}, {13'sd2678, 13'sd2645, 11'sd987}},
{{11'sd-653, 10'sd-479, 13'sd-2245}, {12'sd1475, 13'sd2859, 13'sd-2352}, {12'sd-1821, 13'sd2096, 12'sd-1300}},
{{13'sd-3070, 12'sd1030, 11'sd941}, {13'sd3038, 9'sd-209, 12'sd1698}, {8'sd-91, 12'sd1197, 13'sd2478}},
{{14'sd4647, 12'sd-1289, 14'sd4202}, {12'sd1697, 12'sd-2043, 13'sd2244}, {13'sd2077, 13'sd-2289, 10'sd-418}},
{{12'sd-1563, 13'sd-2485, 7'sd60}, {12'sd1301, 13'sd2789, 12'sd1292}, {13'sd-2214, 11'sd606, 12'sd-1209}},
{{9'sd-192, 12'sd1270, 12'sd-1459}, {13'sd-2322, 12'sd1507, 10'sd482}, {12'sd1824, 12'sd1457, 10'sd-353}},
{{12'sd-1651, 9'sd-211, 9'sd140}, {12'sd1449, 13'sd2459, 12'sd1603}, {10'sd-273, 11'sd-730, 12'sd1287}},
{{12'sd1247, 10'sd391, 11'sd804}, {10'sd-507, 10'sd373, 13'sd-2500}, {9'sd-173, 13'sd-2177, 13'sd-2384}},
{{12'sd-1761, 12'sd-1815, 13'sd-3438}, {13'sd2449, 13'sd-3018, 10'sd298}, {9'sd209, 13'sd-3196, 13'sd-3816}},
{{12'sd-1185, 11'sd955, 10'sd-501}, {12'sd1113, 9'sd-136, 9'sd144}, {12'sd1148, 12'sd1873, 13'sd-2552}},
{{13'sd2079, 13'sd3343, 9'sd-185}, {10'sd-384, 10'sd-306, 9'sd-208}, {11'sd-551, 11'sd-1000, 11'sd933}},
{{12'sd-1978, 10'sd313, 11'sd885}, {12'sd-1886, 12'sd1870, 12'sd1384}, {10'sd472, 9'sd-212, 11'sd-602}},
{{12'sd1627, 11'sd707, 12'sd-1836}, {13'sd2485, 13'sd2870, 12'sd-1648}, {10'sd-306, 12'sd-1311, 12'sd2006}},
{{11'sd777, 10'sd356, 13'sd-2776}, {11'sd599, 13'sd3103, 12'sd-1660}, {11'sd871, 11'sd861, 11'sd571}},
{{12'sd1276, 12'sd1570, 10'sd467}, {12'sd-1831, 11'sd612, 11'sd995}, {13'sd2889, 11'sd807, 11'sd-539}},
{{11'sd779, 12'sd2008, 8'sd105}, {10'sd-431, 12'sd2042, 12'sd-2034}, {11'sd956, 9'sd-173, 11'sd-623}},
{{12'sd-1101, 13'sd-2711, 12'sd-1961}, {11'sd852, 11'sd-924, 12'sd-1055}, {12'sd-1468, 13'sd-3247, 13'sd-2404}},
{{12'sd-1066, 13'sd3289, 11'sd-548}, {13'sd-2054, 13'sd-2600, 10'sd401}, {13'sd-2724, 11'sd-996, 11'sd-705}},
{{13'sd3218, 12'sd1326, 13'sd2101}, {11'sd1002, 13'sd-2332, 12'sd-1407}, {13'sd-2628, 12'sd1707, 11'sd699}},
{{13'sd-2809, 12'sd-1826, 13'sd-2695}, {11'sd-826, 7'sd-45, 11'sd-537}, {13'sd2973, 13'sd-2081, 12'sd1465}},
{{9'sd-198, 12'sd-1817, 12'sd1633}, {13'sd2504, 11'sd983, 12'sd2016}, {12'sd-1821, 13'sd2048, 11'sd-515}},
{{12'sd-1908, 12'sd1299, 8'sd89}, {13'sd2128, 12'sd-1157, 12'sd-1087}, {12'sd1416, 11'sd595, 13'sd-2088}},
{{12'sd-1557, 12'sd1097, 12'sd-1200}, {11'sd-900, 12'sd-1081, 12'sd-1939}, {5'sd12, 10'sd449, 11'sd-1013}},
{{12'sd1643, 9'sd-200, 10'sd-305}, {13'sd3159, 12'sd-1037, 13'sd-2155}, {12'sd1127, 13'sd3447, 12'sd1660}},
{{12'sd1058, 12'sd1579, 8'sd-119}, {9'sd234, 13'sd2259, 8'sd109}, {12'sd-1303, 12'sd-1381, 12'sd1553}},
{{13'sd2476, 12'sd-1573, 12'sd-1770}, {8'sd-104, 9'sd-157, 12'sd1883}, {13'sd2958, 12'sd-1496, 9'sd-235}},
{{10'sd-392, 11'sd642, 14'sd-4281}, {11'sd-667, 11'sd643, 10'sd309}, {12'sd1806, 12'sd-1279, 12'sd-1417}},
{{11'sd-667, 13'sd2296, 12'sd1048}, {13'sd-2412, 10'sd-348, 12'sd-1703}, {11'sd674, 10'sd361, 11'sd526}},
{{13'sd2396, 13'sd2323, 9'sd-162}, {11'sd-605, 10'sd-355, 13'sd-2128}, {12'sd-1407, 13'sd2118, 11'sd-742}},
{{13'sd-3446, 13'sd2651, 11'sd-669}, {11'sd729, 11'sd880, 12'sd-1046}, {13'sd-2209, 12'sd1927, 12'sd-1394}},
{{11'sd-907, 11'sd-633, 11'sd-560}, {11'sd730, 13'sd3027, 7'sd61}, {11'sd-546, 11'sd564, 12'sd-1576}},
{{13'sd2219, 13'sd-2227, 11'sd560}, {11'sd776, 9'sd189, 12'sd-1026}, {8'sd119, 11'sd-621, 6'sd29}},
{{12'sd-1129, 12'sd1565, 10'sd361}, {12'sd-1244, 13'sd2723, 11'sd961}, {10'sd345, 10'sd-362, 10'sd-470}},
{{10'sd-280, 12'sd-1381, 10'sd-346}, {11'sd557, 12'sd-1907, 13'sd-2373}, {12'sd1876, 11'sd759, 12'sd-1864}},
{{11'sd686, 10'sd-450, 12'sd-1723}, {10'sd-497, 12'sd1616, 11'sd800}, {12'sd1786, 13'sd-2503, 9'sd-253}},
{{11'sd-781, 12'sd1243, 11'sd821}, {11'sd-539, 12'sd-1425, 11'sd1004}, {9'sd-245, 10'sd257, 11'sd796}},
{{12'sd-1770, 11'sd-586, 8'sd-72}, {14'sd-4301, 13'sd2056, 13'sd2355}, {13'sd-3047, 12'sd-1893, 12'sd-1154}},
{{12'sd1066, 12'sd-1601, 10'sd-434}, {12'sd-1164, 13'sd-2547, 9'sd161}, {12'sd-1491, 12'sd1448, 10'sd-464}},
{{12'sd1265, 8'sd-125, 13'sd-2742}, {6'sd27, 13'sd-2662, 12'sd-1360}, {11'sd707, 12'sd-1426, 10'sd-384}},
{{13'sd-2407, 11'sd-634, 12'sd-1714}, {11'sd-1009, 9'sd223, 11'sd521}, {12'sd-1999, 12'sd-1662, 12'sd-1364}},
{{11'sd805, 11'sd856, 13'sd2462}, {12'sd-1145, 11'sd-539, 11'sd628}, {13'sd-3665, 11'sd738, 11'sd986}},
{{12'sd-1926, 12'sd1848, 7'sd-49}, {11'sd-908, 12'sd1384, 12'sd1701}, {11'sd-991, 13'sd-2998, 11'sd-871}},
{{12'sd-1245, 12'sd1943, 10'sd416}, {12'sd-1788, 12'sd-1418, 9'sd189}, {11'sd774, 12'sd-1121, 12'sd1463}},
{{13'sd-2725, 12'sd-1966, 14'sd-4259}, {14'sd-5592, 13'sd-3285, 12'sd1287}, {12'sd-1558, 14'sd-4509, 11'sd-835}},
{{12'sd1424, 11'sd-706, 10'sd-401}, {12'sd1610, 13'sd3296, 6'sd17}, {12'sd-1957, 13'sd2731, 12'sd-1816}},
{{9'sd177, 12'sd1379, 10'sd380}, {12'sd-1508, 11'sd993, 13'sd-2448}, {11'sd952, 11'sd-783, 12'sd1325}},
{{11'sd766, 10'sd378, 11'sd-711}, {13'sd2529, 13'sd-2558, 10'sd-494}, {4'sd-7, 13'sd-3595, 11'sd-853}},
{{10'sd-455, 12'sd1632, 11'sd864}, {12'sd-1595, 9'sd200, 12'sd-1147}, {7'sd-53, 10'sd-476, 12'sd1176}},
{{13'sd2435, 12'sd1385, 12'sd-1136}, {12'sd1300, 13'sd2705, 12'sd2036}, {11'sd934, 13'sd2365, 11'sd-530}},
{{9'sd-148, 12'sd-1578, 12'sd1270}, {12'sd1461, 12'sd-1259, 12'sd1623}, {12'sd1377, 11'sd715, 11'sd515}},
{{12'sd-1578, 10'sd-493, 13'sd3431}, {12'sd1209, 9'sd-183, 10'sd404}, {12'sd1680, 10'sd-290, 10'sd419}},
{{12'sd1326, 12'sd-1768, 10'sd-367}, {11'sd-539, 8'sd74, 11'sd-662}, {12'sd-1192, 12'sd1909, 12'sd1582}},
{{12'sd2016, 13'sd2122, 10'sd261}, {10'sd-306, 12'sd-1126, 12'sd1094}, {12'sd-1349, 12'sd-1090, 12'sd1125}},
{{12'sd1205, 13'sd-2449, 10'sd-383}, {13'sd2572, 13'sd-2342, 11'sd-994}, {13'sd2929, 12'sd-1446, 13'sd-3728}},
{{12'sd-1771, 11'sd881, 12'sd-1890}, {12'sd-1213, 10'sd372, 12'sd1138}, {13'sd2348, 9'sd-240, 12'sd-1869}},
{{12'sd1031, 12'sd-1397, 13'sd-2165}, {4'sd-5, 12'sd1434, 13'sd2273}, {12'sd-1540, 9'sd227, 9'sd-164}},
{{12'sd-1821, 11'sd-845, 11'sd-850}, {12'sd1143, 13'sd2322, 12'sd1458}, {13'sd2122, 11'sd-757, 13'sd2756}},
{{11'sd-973, 11'sd-568, 12'sd-1506}, {11'sd-591, 13'sd2287, 11'sd-902}, {12'sd1615, 11'sd-732, 13'sd2130}},
{{11'sd-561, 11'sd858, 12'sd-2016}, {13'sd2062, 10'sd-397, 13'sd-2612}, {12'sd1589, 13'sd-2405, 13'sd-2346}},
{{11'sd654, 12'sd-1209, 13'sd3443}, {11'sd795, 10'sd-437, 10'sd280}, {11'sd-635, 11'sd868, 13'sd-2395}}},
{
{{12'sd-1300, 11'sd649, 9'sd-254}, {9'sd230, 11'sd-771, 13'sd-2193}, {10'sd496, 11'sd893, 12'sd-1507}},
{{13'sd2504, 13'sd-2094, 13'sd2232}, {12'sd-1384, 13'sd2727, 11'sd-992}, {10'sd-306, 8'sd-120, 12'sd1926}},
{{13'sd3118, 13'sd-2163, 11'sd796}, {12'sd-1764, 13'sd-2735, 11'sd894}, {11'sd914, 12'sd1099, 13'sd-3552}},
{{11'sd-686, 12'sd1192, 13'sd3009}, {13'sd3087, 13'sd2805, 13'sd2172}, {13'sd-2197, 12'sd-1730, 12'sd-1233}},
{{10'sd368, 11'sd946, 13'sd2431}, {11'sd-556, 12'sd-1190, 10'sd275}, {12'sd-1526, 12'sd1489, 12'sd-1805}},
{{13'sd-2602, 13'sd2289, 9'sd136}, {9'sd174, 12'sd1888, 10'sd-269}, {11'sd-580, 13'sd2414, 12'sd1067}},
{{11'sd-662, 10'sd339, 11'sd-722}, {12'sd1296, 13'sd-2278, 11'sd-587}, {13'sd3253, 11'sd898, 12'sd1176}},
{{12'sd-1940, 13'sd2792, 12'sd1449}, {13'sd2777, 9'sd-213, 10'sd-510}, {12'sd-1367, 8'sd-81, 11'sd-793}},
{{12'sd1411, 12'sd-2005, 12'sd-1241}, {12'sd-1044, 8'sd108, 13'sd-2097}, {13'sd-3176, 12'sd1556, 12'sd-1554}},
{{12'sd1155, 13'sd-2461, 11'sd-793}, {13'sd-2611, 7'sd33, 12'sd-1273}, {12'sd1655, 11'sd836, 12'sd1592}},
{{13'sd2272, 13'sd2334, 10'sd333}, {12'sd1567, 12'sd-1362, 12'sd1685}, {12'sd-1433, 10'sd394, 13'sd-2411}},
{{12'sd-1219, 13'sd-2112, 13'sd2699}, {11'sd-1015, 11'sd940, 12'sd1683}, {10'sd355, 12'sd-1573, 10'sd-394}},
{{13'sd-3466, 12'sd-1608, 12'sd-1147}, {12'sd1428, 12'sd-1650, 12'sd-2028}, {12'sd-1041, 10'sd395, 11'sd-880}},
{{12'sd1542, 13'sd-2770, 13'sd2528}, {6'sd21, 10'sd-483, 10'sd-416}, {11'sd863, 13'sd-2309, 12'sd1358}},
{{11'sd625, 12'sd1645, 11'sd895}, {12'sd-1807, 12'sd-1245, 12'sd-1310}, {13'sd-2385, 12'sd1212, 11'sd855}},
{{10'sd332, 11'sd1015, 13'sd-2099}, {13'sd2198, 12'sd1566, 13'sd2090}, {9'sd-154, 11'sd-886, 11'sd531}},
{{13'sd-2249, 13'sd-2344, 9'sd193}, {13'sd-2067, 9'sd-143, 13'sd2322}, {12'sd-2035, 12'sd1561, 12'sd-2021}},
{{12'sd1779, 10'sd510, 12'sd1038}, {12'sd-1311, 11'sd753, 11'sd643}, {12'sd-1416, 10'sd-396, 12'sd1812}},
{{13'sd2782, 12'sd-1373, 12'sd-1461}, {11'sd-694, 12'sd1151, 12'sd1709}, {12'sd-1344, 13'sd2498, 11'sd-1015}},
{{11'sd-777, 12'sd-1470, 11'sd522}, {12'sd-1315, 12'sd-1834, 13'sd-2138}, {12'sd1535, 10'sd-278, 13'sd2425}},
{{9'sd233, 12'sd-1363, 11'sd-915}, {11'sd841, 12'sd-2026, 11'sd-687}, {12'sd-2042, 12'sd-1803, 11'sd-721}},
{{12'sd-1427, 13'sd3027, 11'sd608}, {10'sd-265, 13'sd-2446, 12'sd1182}, {13'sd-2438, 11'sd-1015, 12'sd-1546}},
{{13'sd2554, 9'sd249, 12'sd1156}, {13'sd-2577, 12'sd1617, 8'sd90}, {13'sd-2083, 11'sd-571, 13'sd-2632}},
{{12'sd-1058, 13'sd2378, 11'sd-717}, {12'sd1354, 11'sd721, 11'sd-534}, {10'sd-486, 12'sd-1640, 11'sd-782}},
{{12'sd-1890, 10'sd459, 12'sd-1444}, {11'sd764, 10'sd266, 12'sd1600}, {11'sd957, 13'sd2665, 11'sd953}},
{{11'sd592, 9'sd-160, 13'sd2668}, {10'sd-509, 10'sd-340, 11'sd696}, {13'sd2367, 13'sd2487, 10'sd-394}},
{{12'sd1616, 12'sd1403, 11'sd530}, {13'sd2160, 12'sd1157, 10'sd-304}, {13'sd2395, 13'sd-2704, 13'sd2469}},
{{12'sd1100, 12'sd1338, 12'sd1602}, {13'sd3203, 13'sd-2216, 12'sd-1517}, {12'sd1377, 13'sd3476, 13'sd2317}},
{{10'sd406, 13'sd2305, 11'sd639}, {10'sd495, 12'sd1085, 13'sd-2212}, {13'sd-2066, 13'sd-2893, 13'sd2052}},
{{12'sd2041, 10'sd370, 11'sd-537}, {12'sd-1451, 8'sd-69, 8'sd66}, {12'sd1382, 12'sd2009, 13'sd2088}},
{{10'sd386, 4'sd-5, 13'sd-2228}, {12'sd-1179, 13'sd2326, 12'sd-1842}, {13'sd3195, 13'sd2621, 13'sd2480}},
{{12'sd1045, 11'sd-878, 13'sd2219}, {12'sd1265, 12'sd-1791, 12'sd1518}, {11'sd-901, 12'sd-2028, 11'sd703}},
{{13'sd2488, 12'sd1042, 12'sd-1597}, {13'sd-2113, 12'sd1468, 13'sd-3248}, {13'sd2646, 12'sd1082, 12'sd1969}},
{{11'sd956, 12'sd-1622, 13'sd2277}, {11'sd774, 10'sd-315, 13'sd2348}, {12'sd1852, 12'sd-1331, 9'sd-130}},
{{9'sd205, 12'sd-1263, 13'sd2111}, {12'sd-1530, 13'sd2423, 10'sd315}, {12'sd1210, 12'sd-2038, 13'sd-2409}},
{{9'sd-131, 8'sd100, 12'sd-1393}, {12'sd1950, 10'sd-495, 12'sd1141}, {13'sd-2949, 12'sd1466, 11'sd-550}},
{{12'sd1779, 13'sd-2180, 11'sd-525}, {12'sd-1711, 11'sd-715, 11'sd-733}, {12'sd-1164, 13'sd2697, 12'sd-1734}},
{{13'sd2743, 11'sd538, 13'sd-2183}, {11'sd805, 13'sd2442, 13'sd2661}, {12'sd1281, 12'sd1369, 13'sd-2564}},
{{13'sd2690, 10'sd380, 13'sd2636}, {12'sd1713, 7'sd-56, 11'sd783}, {12'sd1571, 11'sd-677, 12'sd1191}},
{{13'sd2117, 9'sd-223, 10'sd330}, {11'sd529, 13'sd2317, 11'sd721}, {10'sd328, 13'sd2213, 12'sd1091}},
{{11'sd-740, 12'sd-1409, 12'sd-1439}, {12'sd-1223, 12'sd-1257, 11'sd-963}, {11'sd-659, 12'sd1095, 11'sd532}},
{{13'sd-2590, 12'sd1138, 11'sd583}, {12'sd1646, 11'sd-882, 9'sd136}, {10'sd-487, 12'sd-1978, 13'sd-2867}},
{{8'sd82, 13'sd-2769, 11'sd-927}, {7'sd37, 9'sd-221, 12'sd1666}, {11'sd-825, 12'sd1893, 11'sd900}},
{{12'sd-1635, 12'sd-1083, 8'sd117}, {12'sd-1545, 11'sd-557, 12'sd-1211}, {13'sd-2468, 13'sd-2731, 12'sd-1130}},
{{12'sd-1867, 12'sd-2015, 12'sd-1323}, {12'sd1748, 12'sd-1395, 12'sd-1353}, {12'sd1313, 12'sd1590, 13'sd-2584}},
{{11'sd-779, 12'sd1177, 9'sd213}, {11'sd668, 13'sd2729, 12'sd2022}, {11'sd899, 11'sd-614, 13'sd2284}},
{{13'sd-2538, 13'sd2602, 9'sd224}, {13'sd-2325, 13'sd-2355, 12'sd-1216}, {12'sd1085, 13'sd-2527, 9'sd208}},
{{13'sd-2764, 10'sd-496, 11'sd1019}, {12'sd-1679, 12'sd-1401, 12'sd-1984}, {8'sd-112, 12'sd-1936, 13'sd-3120}},
{{13'sd2542, 9'sd133, 6'sd-26}, {9'sd-225, 12'sd-1459, 13'sd-2085}, {11'sd-622, 11'sd555, 11'sd813}},
{{11'sd766, 12'sd1350, 12'sd1972}, {8'sd119, 12'sd1275, 12'sd-1722}, {12'sd1725, 12'sd-1389, 12'sd1919}},
{{13'sd-2133, 9'sd-143, 9'sd249}, {10'sd354, 9'sd182, 4'sd6}, {13'sd-2605, 11'sd-524, 10'sd-427}},
{{12'sd1956, 9'sd184, 8'sd111}, {9'sd-150, 13'sd-2647, 12'sd1419}, {13'sd-2336, 11'sd640, 13'sd2255}},
{{13'sd-2331, 13'sd2340, 13'sd2607}, {13'sd-2548, 12'sd-1458, 13'sd2292}, {11'sd-566, 13'sd2413, 12'sd-1092}},
{{8'sd127, 13'sd-2681, 11'sd-711}, {13'sd2656, 11'sd-898, 12'sd-1407}, {13'sd2362, 11'sd-873, 10'sd269}},
{{13'sd3089, 13'sd2282, 9'sd-210}, {12'sd1245, 12'sd1054, 11'sd-751}, {7'sd62, 9'sd-146, 13'sd-2299}},
{{13'sd-2991, 10'sd385, 12'sd1915}, {12'sd1679, 12'sd1441, 11'sd-798}, {13'sd-2289, 11'sd-671, 13'sd-2304}},
{{12'sd-1522, 11'sd863, 12'sd2027}, {12'sd-1872, 8'sd-77, 13'sd2167}, {10'sd-431, 11'sd637, 12'sd1467}},
{{13'sd-2052, 11'sd1010, 11'sd-742}, {11'sd830, 9'sd-181, 12'sd1148}, {13'sd2107, 9'sd129, 12'sd-1485}},
{{13'sd-2065, 12'sd-1311, 9'sd-185}, {12'sd-1054, 12'sd-1252, 11'sd658}, {13'sd3484, 12'sd-1697, 12'sd-1102}},
{{13'sd-3235, 3'sd3, 12'sd1239}, {13'sd-2359, 12'sd-1304, 12'sd-1624}, {9'sd207, 11'sd953, 12'sd-1529}},
{{10'sd-322, 13'sd-2630, 12'sd1543}, {12'sd-1839, 13'sd2056, 12'sd1666}, {12'sd-1535, 12'sd-1897, 11'sd841}},
{{10'sd-380, 9'sd239, 12'sd-1367}, {11'sd-848, 11'sd618, 13'sd2705}, {12'sd-1510, 12'sd-1955, 12'sd-1987}},
{{13'sd2396, 12'sd1964, 11'sd-800}, {10'sd412, 12'sd-1698, 13'sd-2623}, {13'sd-3113, 13'sd-2803, 12'sd1521}},
{{12'sd1095, 12'sd1998, 12'sd-1185}, {13'sd2668, 12'sd-1839, 10'sd335}, {12'sd-1148, 12'sd1746, 13'sd-2995}}},
{
{{12'sd1155, 12'sd-1419, 13'sd-3048}, {13'sd2191, 10'sd-264, 12'sd1068}, {11'sd929, 13'sd2086, 13'sd2223}},
{{11'sd-940, 13'sd-2725, 12'sd1937}, {12'sd-1575, 12'sd1346, 8'sd99}, {12'sd1862, 12'sd1097, 12'sd1586}},
{{11'sd1002, 13'sd-3470, 13'sd-3070}, {13'sd-3057, 11'sd728, 13'sd2287}, {10'sd464, 12'sd1948, 12'sd1680}},
{{13'sd2711, 12'sd1080, 11'sd-846}, {10'sd-283, 11'sd519, 12'sd1236}, {13'sd2772, 12'sd1722, 8'sd-126}},
{{12'sd-1459, 9'sd130, 12'sd1981}, {12'sd1837, 11'sd-766, 11'sd521}, {13'sd-2422, 12'sd1409, 13'sd-2141}},
{{10'sd-305, 12'sd-1093, 12'sd-1390}, {10'sd440, 11'sd1002, 12'sd1809}, {12'sd-2018, 12'sd-1764, 10'sd-495}},
{{9'sd-211, 8'sd108, 7'sd52}, {12'sd1866, 11'sd-631, 11'sd985}, {9'sd137, 12'sd-1080, 12'sd-1411}},
{{12'sd-1592, 12'sd-1887, 11'sd-908}, {11'sd660, 9'sd-152, 13'sd-2445}, {12'sd-1904, 13'sd2338, 12'sd1410}},
{{11'sd569, 12'sd-1672, 11'sd-534}, {13'sd2465, 13'sd2256, 12'sd1076}, {13'sd-2523, 10'sd-268, 12'sd-1780}},
{{12'sd-1299, 13'sd2071, 12'sd1952}, {12'sd-1964, 7'sd-34, 12'sd1665}, {13'sd-2565, 13'sd-2230, 12'sd-1687}},
{{13'sd3219, 13'sd3239, 11'sd575}, {12'sd-1201, 13'sd2339, 12'sd1428}, {10'sd319, 12'sd1573, 11'sd-662}},
{{11'sd-618, 13'sd2397, 12'sd1757}, {13'sd-2507, 13'sd-2384, 10'sd-277}, {11'sd531, 11'sd590, 12'sd1899}},
{{12'sd1642, 13'sd3156, 10'sd338}, {12'sd-1427, 11'sd867, 11'sd536}, {13'sd-2529, 12'sd-1217, 12'sd-2043}},
{{9'sd-215, 13'sd-2411, 12'sd1274}, {11'sd-799, 13'sd-2755, 12'sd-1995}, {12'sd-1345, 10'sd-397, 13'sd-2322}},
{{12'sd1924, 13'sd-2584, 12'sd-1490}, {7'sd-54, 13'sd-2415, 12'sd-1462}, {12'sd-1309, 11'sd1023, 12'sd1440}},
{{12'sd1922, 11'sd691, 12'sd-1029}, {13'sd2848, 12'sd1118, 11'sd604}, {12'sd1453, 12'sd1829, 11'sd-525}},
{{13'sd-2779, 13'sd-2264, 10'sd-463}, {12'sd-1714, 9'sd-182, 12'sd-1633}, {11'sd-568, 11'sd519, 13'sd-2416}},
{{11'sd-521, 12'sd-2023, 12'sd1799}, {10'sd365, 13'sd-2358, 11'sd-648}, {11'sd-834, 8'sd71, 13'sd2338}},
{{13'sd2426, 13'sd2191, 13'sd2587}, {9'sd165, 11'sd968, 12'sd-1827}, {12'sd-1605, 12'sd1681, 12'sd1151}},
{{13'sd2999, 12'sd1740, 13'sd3094}, {12'sd-1747, 12'sd-1936, 10'sd408}, {12'sd1146, 13'sd-2071, 12'sd-1058}},
{{12'sd-1380, 8'sd-122, 13'sd-2287}, {13'sd-2828, 12'sd1045, 13'sd-2220}, {13'sd-2095, 13'sd2696, 12'sd-1540}},
{{12'sd1467, 12'sd1794, 12'sd-1337}, {12'sd1094, 12'sd1592, 12'sd-1335}, {12'sd1128, 12'sd-1208, 11'sd838}},
{{11'sd-953, 12'sd1868, 10'sd298}, {8'sd73, 8'sd-121, 9'sd-212}, {12'sd-1159, 12'sd1073, 10'sd280}},
{{13'sd2497, 13'sd-2518, 12'sd1932}, {8'sd-106, 8'sd69, 12'sd-1300}, {13'sd2399, 12'sd-1902, 12'sd1687}},
{{11'sd828, 12'sd1176, 11'sd-552}, {8'sd-92, 12'sd-1500, 11'sd895}, {11'sd-889, 13'sd2897, 10'sd-346}},
{{12'sd1639, 12'sd-1335, 11'sd-580}, {12'sd-1659, 11'sd-839, 8'sd-70}, {13'sd2649, 11'sd-514, 10'sd298}},
{{12'sd-1605, 11'sd792, 12'sd1723}, {13'sd-2577, 11'sd732, 12'sd-1772}, {13'sd2291, 12'sd-1141, 12'sd1697}},
{{12'sd-1194, 13'sd-2692, 12'sd1274}, {8'sd76, 12'sd-1819, 10'sd277}, {11'sd-670, 13'sd-3253, 12'sd1711}},
{{11'sd-743, 12'sd1900, 12'sd-1781}, {13'sd2460, 12'sd-1373, 12'sd-1792}, {13'sd-2093, 12'sd1592, 10'sd-303}},
{{13'sd-2205, 12'sd1906, 12'sd1967}, {12'sd1829, 13'sd2166, 12'sd1830}, {12'sd-1329, 9'sd184, 10'sd443}},
{{11'sd632, 12'sd1403, 13'sd2628}, {12'sd-1697, 4'sd-7, 7'sd35}, {10'sd-437, 13'sd-2341, 10'sd479}},
{{13'sd-2882, 9'sd193, 13'sd-3265}, {12'sd-1195, 12'sd1498, 6'sd19}, {13'sd-2576, 12'sd1563, 12'sd1763}},
{{11'sd-915, 12'sd1621, 12'sd-1948}, {11'sd-766, 10'sd401, 11'sd-953}, {13'sd2452, 11'sd747, 12'sd1275}},
{{12'sd1737, 13'sd-2569, 11'sd-929}, {13'sd2161, 12'sd-1749, 11'sd-548}, {12'sd1304, 12'sd-1346, 12'sd1560}},
{{11'sd-635, 12'sd-1335, 13'sd-2184}, {13'sd-2051, 11'sd955, 12'sd-1853}, {12'sd-1253, 12'sd1719, 12'sd1539}},
{{10'sd496, 13'sd-2188, 12'sd1140}, {12'sd1901, 13'sd-2192, 12'sd1580}, {12'sd1074, 12'sd2023, 12'sd-1270}},
{{9'sd-212, 12'sd-1716, 12'sd2032}, {12'sd-1853, 12'sd-1509, 13'sd2907}, {12'sd1900, 10'sd460, 12'sd-1958}},
{{13'sd-2233, 13'sd2366, 12'sd1881}, {11'sd779, 12'sd-1775, 10'sd-380}, {13'sd2507, 12'sd1755, 13'sd2310}},
{{13'sd-2283, 12'sd1309, 12'sd1394}, {13'sd2194, 12'sd1407, 11'sd-712}, {13'sd2576, 12'sd-1798, 11'sd-685}},
{{12'sd-1094, 11'sd-700, 10'sd367}, {10'sd414, 11'sd-979, 12'sd-1082}, {13'sd2116, 12'sd-1791, 13'sd2713}},
{{12'sd1587, 12'sd1849, 13'sd3404}, {12'sd-1272, 11'sd616, 13'sd2318}, {12'sd1593, 12'sd-1346, 12'sd2009}},
{{12'sd1550, 12'sd-1415, 12'sd-1860}, {10'sd462, 13'sd2404, 12'sd-1387}, {8'sd65, 11'sd803, 10'sd-316}},
{{12'sd1890, 12'sd1765, 12'sd1700}, {12'sd-1394, 9'sd-236, 10'sd-340}, {12'sd-1280, 13'sd2861, 12'sd-1828}},
{{13'sd2836, 11'sd1018, 12'sd-1880}, {13'sd2843, 12'sd1430, 13'sd2871}, {13'sd2170, 12'sd1791, 12'sd-1952}},
{{13'sd-2140, 12'sd1646, 12'sd1547}, {9'sd-160, 12'sd-1268, 13'sd2746}, {10'sd350, 12'sd1409, 12'sd-1281}},
{{13'sd2051, 8'sd74, 12'sd-1765}, {12'sd-1885, 12'sd1111, 9'sd232}, {10'sd367, 9'sd170, 12'sd1811}},
{{12'sd1851, 10'sd-422, 12'sd1978}, {10'sd-345, 11'sd-919, 12'sd-1827}, {12'sd1065, 12'sd1504, 11'sd803}},
{{11'sd888, 12'sd-1729, 12'sd-1042}, {13'sd2652, 10'sd471, 12'sd1920}, {11'sd924, 13'sd-2052, 11'sd756}},
{{11'sd-905, 12'sd-1773, 9'sd-242}, {10'sd-502, 12'sd1826, 13'sd-2197}, {12'sd-1808, 11'sd-568, 12'sd1270}},
{{10'sd419, 13'sd2307, 12'sd1699}, {13'sd2732, 12'sd-1229, 10'sd-495}, {13'sd-2424, 7'sd-41, 12'sd-1901}},
{{13'sd2790, 11'sd-884, 13'sd-2604}, {13'sd2317, 13'sd-2101, 11'sd-631}, {10'sd-295, 12'sd-1728, 13'sd-3047}},
{{12'sd1788, 11'sd832, 9'sd138}, {10'sd406, 12'sd-1057, 13'sd2377}, {7'sd33, 12'sd-1868, 11'sd915}},
{{12'sd1820, 2'sd1, 11'sd626}, {12'sd1241, 10'sd409, 11'sd840}, {12'sd-1923, 9'sd-243, 12'sd-1141}},
{{12'sd-1651, 10'sd322, 11'sd612}, {12'sd-1456, 7'sd41, 10'sd380}, {11'sd905, 11'sd880, 13'sd2403}},
{{13'sd2446, 13'sd2532, 10'sd-271}, {8'sd-65, 11'sd-884, 12'sd-1224}, {11'sd-594, 13'sd-2375, 10'sd257}},
{{12'sd-1812, 12'sd-1955, 11'sd-578}, {11'sd-674, 12'sd-1473, 13'sd-2262}, {8'sd-115, 13'sd-2418, 13'sd2278}},
{{13'sd2543, 12'sd-1821, 12'sd1834}, {12'sd-1333, 6'sd30, 11'sd574}, {10'sd-258, 12'sd1686, 12'sd1124}},
{{11'sd707, 13'sd2392, 10'sd-271}, {12'sd-1606, 9'sd177, 13'sd-2320}, {13'sd-2281, 10'sd353, 13'sd2707}},
{{9'sd174, 11'sd980, 10'sd458}, {8'sd101, 8'sd-80, 11'sd-573}, {11'sd818, 13'sd2471, 13'sd-2094}},
{{13'sd-2433, 13'sd-2544, 13'sd-2990}, {12'sd1728, 13'sd2319, 12'sd1777}, {12'sd-1842, 11'sd884, 13'sd-2168}},
{{11'sd671, 9'sd-155, 13'sd2269}, {13'sd-2564, 12'sd-1959, 12'sd1166}, {10'sd-267, 12'sd-1613, 13'sd-2755}},
{{12'sd-1862, 8'sd83, 12'sd-1520}, {13'sd-2545, 13'sd2158, 11'sd-906}, {12'sd1603, 12'sd1180, 12'sd-1929}},
{{13'sd2578, 11'sd-532, 10'sd345}, {12'sd1353, 12'sd1769, 11'sd1014}, {13'sd2601, 9'sd148, 12'sd1588}},
{{12'sd-1643, 12'sd-1717, 13'sd-2605}, {12'sd-1261, 12'sd-1436, 11'sd-531}, {13'sd-2327, 12'sd1123, 10'sd-389}}},
{
{{10'sd-481, 13'sd2350, 12'sd-1644}, {13'sd2176, 12'sd-1675, 6'sd17}, {10'sd-501, 12'sd-1325, 12'sd1364}},
{{12'sd1358, 12'sd1782, 13'sd2223}, {9'sd242, 13'sd2303, 13'sd-2962}, {11'sd555, 12'sd-1357, 10'sd452}},
{{12'sd-1294, 11'sd579, 13'sd2245}, {11'sd-736, 12'sd-1933, 11'sd909}, {14'sd-4726, 13'sd-3981, 13'sd-2801}},
{{12'sd-1957, 10'sd-332, 9'sd-183}, {12'sd-1307, 10'sd-423, 13'sd2194}, {11'sd-917, 13'sd-2650, 11'sd772}},
{{10'sd-501, 13'sd-3131, 13'sd2179}, {12'sd-1853, 8'sd69, 13'sd2416}, {12'sd1389, 11'sd-761, 12'sd1602}},
{{12'sd1722, 11'sd710, 9'sd137}, {7'sd39, 13'sd-2840, 10'sd350}, {12'sd-1203, 13'sd2366, 12'sd-1073}},
{{12'sd-1137, 13'sd-3098, 13'sd-2790}, {12'sd1162, 12'sd1647, 12'sd-1055}, {9'sd199, 12'sd-1029, 12'sd1686}},
{{12'sd1549, 12'sd1160, 11'sd-547}, {12'sd-1398, 11'sd691, 13'sd-2163}, {12'sd1416, 11'sd771, 13'sd2149}},
{{13'sd-2530, 9'sd244, 13'sd2382}, {13'sd2540, 12'sd-1361, 12'sd-1182}, {12'sd1412, 13'sd-2340, 12'sd1280}},
{{11'sd665, 13'sd-2078, 12'sd1857}, {10'sd296, 12'sd1509, 13'sd-2502}, {13'sd2527, 11'sd-556, 11'sd810}},
{{13'sd-2823, 12'sd-1586, 12'sd-1726}, {6'sd17, 12'sd-1722, 12'sd-1410}, {13'sd-2191, 9'sd197, 13'sd2269}},
{{12'sd-1404, 13'sd2268, 12'sd1882}, {10'sd441, 12'sd-1461, 13'sd-2071}, {12'sd-1466, 10'sd-268, 13'sd-2405}},
{{12'sd-1309, 11'sd761, 12'sd1387}, {13'sd2184, 7'sd-61, 8'sd-115}, {10'sd257, 12'sd1472, 13'sd2334}},
{{9'sd-213, 11'sd929, 13'sd2597}, {13'sd2992, 13'sd-2165, 12'sd-1153}, {9'sd-191, 12'sd-1279, 11'sd-662}},
{{10'sd300, 11'sd-901, 12'sd2039}, {12'sd1274, 12'sd1642, 12'sd-1543}, {12'sd1896, 12'sd1901, 12'sd-1089}},
{{11'sd-522, 13'sd2445, 10'sd-485}, {10'sd-484, 11'sd679, 12'sd1877}, {12'sd1129, 9'sd143, 10'sd-276}},
{{8'sd72, 10'sd375, 11'sd-934}, {12'sd1858, 12'sd1416, 12'sd-1709}, {10'sd-460, 12'sd1998, 12'sd-1356}},
{{10'sd-315, 12'sd1249, 12'sd-1975}, {10'sd492, 11'sd-860, 12'sd1223}, {11'sd1004, 12'sd-2036, 13'sd2341}},
{{12'sd1571, 13'sd2563, 13'sd2400}, {11'sd-545, 12'sd-1606, 13'sd-2288}, {12'sd-1890, 9'sd159, 11'sd-681}},
{{11'sd743, 11'sd824, 9'sd166}, {10'sd-504, 12'sd-1334, 11'sd-1014}, {12'sd1794, 12'sd1991, 12'sd-1639}},
{{12'sd1761, 12'sd1438, 13'sd-2369}, {12'sd1165, 12'sd1947, 9'sd-166}, {9'sd-195, 8'sd-126, 13'sd-3634}},
{{8'sd122, 12'sd-1413, 12'sd-1855}, {12'sd1591, 10'sd-275, 6'sd17}, {13'sd2899, 8'sd66, 10'sd-431}},
{{11'sd946, 12'sd1753, 11'sd-576}, {11'sd-561, 13'sd2141, 12'sd1824}, {13'sd-2528, 12'sd1917, 10'sd-399}},
{{13'sd-2214, 13'sd-2272, 13'sd-2319}, {10'sd299, 13'sd2142, 12'sd1245}, {13'sd-2114, 11'sd-657, 12'sd-1326}},
{{12'sd1241, 12'sd-1835, 9'sd-178}, {13'sd-2422, 13'sd-2059, 13'sd-2191}, {12'sd-1842, 11'sd623, 13'sd2704}},
{{13'sd2192, 12'sd1090, 12'sd-1393}, {12'sd-2036, 11'sd-963, 11'sd772}, {12'sd1939, 13'sd2329, 12'sd1349}},
{{11'sd798, 10'sd360, 12'sd-2000}, {12'sd-1056, 12'sd-1462, 12'sd1210}, {11'sd920, 12'sd-2030, 13'sd2326}},
{{12'sd-1842, 12'sd-1585, 13'sd-2643}, {13'sd2483, 13'sd-2625, 11'sd-796}, {12'sd1285, 12'sd1508, 11'sd-906}},
{{12'sd1626, 8'sd93, 12'sd1909}, {11'sd722, 11'sd-577, 13'sd-2053}, {13'sd2364, 9'sd-148, 13'sd2432}},
{{11'sd-727, 7'sd38, 10'sd-301}, {12'sd1026, 11'sd-994, 12'sd-1209}, {12'sd-1057, 12'sd-1998, 10'sd391}},
{{12'sd-1637, 11'sd-850, 12'sd1321}, {13'sd2808, 11'sd676, 11'sd-939}, {13'sd3164, 11'sd-999, 11'sd786}},
{{11'sd1018, 11'sd-575, 10'sd318}, {13'sd2775, 9'sd254, 13'sd-2599}, {13'sd2752, 11'sd-823, 11'sd-809}},
{{12'sd-1232, 11'sd888, 11'sd-644}, {12'sd1101, 12'sd1752, 12'sd1151}, {11'sd-790, 11'sd584, 13'sd3392}},
{{12'sd-1531, 12'sd-1870, 12'sd-1457}, {10'sd-286, 13'sd3295, 12'sd1261}, {12'sd1574, 13'sd-2429, 11'sd-1009}},
{{12'sd1068, 13'sd2625, 11'sd829}, {11'sd807, 11'sd662, 11'sd948}, {10'sd332, 10'sd370, 11'sd946}},
{{6'sd-17, 12'sd-2003, 11'sd856}, {12'sd-1037, 13'sd2635, 12'sd-1200}, {12'sd1436, 13'sd2146, 13'sd2215}},
{{13'sd-2544, 11'sd514, 12'sd-1657}, {13'sd-2553, 10'sd482, 12'sd-1340}, {12'sd1514, 12'sd1054, 12'sd-1817}},
{{12'sd1292, 12'sd1410, 7'sd45}, {13'sd2936, 11'sd894, 12'sd1490}, {11'sd926, 11'sd981, 12'sd-1177}},
{{11'sd662, 11'sd951, 12'sd1996}, {11'sd923, 13'sd2715, 12'sd-1521}, {12'sd-1988, 10'sd-391, 12'sd1807}},
{{8'sd-107, 10'sd-341, 13'sd-2429}, {11'sd906, 11'sd538, 12'sd1116}, {10'sd-397, 12'sd1714, 10'sd433}},
{{12'sd-1188, 12'sd1671, 14'sd-4125}, {11'sd-843, 13'sd2154, 11'sd-529}, {10'sd-344, 13'sd-2303, 9'sd-242}},
{{13'sd2870, 8'sd97, 12'sd1820}, {11'sd916, 13'sd2209, 11'sd-667}, {10'sd499, 11'sd719, 11'sd-1006}},
{{11'sd712, 12'sd1656, 11'sd634}, {13'sd-2203, 12'sd1938, 12'sd-1051}, {11'sd-520, 12'sd-1189, 13'sd-2613}},
{{10'sd328, 10'sd427, 13'sd2721}, {11'sd-874, 13'sd2317, 13'sd-2236}, {12'sd1122, 13'sd-2143, 10'sd360}},
{{12'sd1149, 12'sd1529, 12'sd1815}, {11'sd-900, 13'sd-3080, 13'sd-2060}, {13'sd-2143, 11'sd-761, 13'sd-2891}},
{{11'sd832, 8'sd-67, 9'sd129}, {12'sd1833, 12'sd-1700, 10'sd-276}, {11'sd525, 12'sd-1480, 13'sd2486}},
{{13'sd-2741, 12'sd-1528, 9'sd-211}, {13'sd2571, 12'sd-1045, 12'sd2027}, {12'sd1583, 12'sd1351, 12'sd-1849}},
{{13'sd2216, 13'sd2244, 12'sd2031}, {13'sd-2599, 12'sd-1273, 12'sd1538}, {11'sd-709, 12'sd-1818, 11'sd-515}},
{{13'sd-2854, 10'sd-284, 12'sd-1231}, {13'sd2463, 12'sd1385, 12'sd1322}, {13'sd-2408, 13'sd2231, 13'sd-2709}},
{{12'sd-1065, 12'sd-1464, 12'sd-1379}, {11'sd944, 13'sd-2555, 12'sd1524}, {14'sd4127, 13'sd3419, 10'sd277}},
{{12'sd-1683, 11'sd-796, 10'sd-459}, {12'sd-1393, 9'sd237, 10'sd382}, {12'sd-1864, 11'sd-619, 12'sd-1616}},
{{13'sd-2809, 9'sd-182, 13'sd-2468}, {9'sd-191, 12'sd-1930, 12'sd1749}, {12'sd-1967, 13'sd-2174, 12'sd-1386}},
{{12'sd1638, 8'sd71, 12'sd-1675}, {12'sd-1773, 13'sd-2669, 13'sd-2658}, {10'sd455, 12'sd1373, 12'sd1555}},
{{6'sd-18, 12'sd-1943, 13'sd-2301}, {9'sd135, 11'sd-843, 12'sd1793}, {11'sd-941, 12'sd-1134, 13'sd-2761}},
{{12'sd1758, 12'sd-1146, 12'sd-1614}, {13'sd2161, 13'sd2141, 12'sd1609}, {11'sd-612, 10'sd-430, 13'sd-3052}},
{{12'sd-1523, 11'sd587, 8'sd-66}, {13'sd-2483, 13'sd-2637, 11'sd-708}, {13'sd-2869, 12'sd-1536, 13'sd2420}},
{{12'sd1768, 10'sd-465, 11'sd-945}, {12'sd-1397, 12'sd-1437, 13'sd-2301}, {13'sd2251, 11'sd882, 12'sd1405}},
{{13'sd3068, 12'sd-1868, 11'sd926}, {10'sd-256, 10'sd-424, 12'sd1906}, {11'sd979, 11'sd1013, 12'sd1958}},
{{11'sd996, 11'sd-694, 12'sd-1362}, {13'sd-2332, 11'sd-716, 12'sd-1862}, {12'sd-1448, 11'sd970, 11'sd-997}},
{{7'sd-60, 12'sd1368, 12'sd-1872}, {12'sd-1579, 13'sd2413, 12'sd-1973}, {13'sd-2652, 11'sd928, 12'sd1323}},
{{12'sd2027, 13'sd-2833, 12'sd1672}, {12'sd1024, 11'sd1019, 11'sd-516}, {11'sd903, 12'sd1225, 11'sd-805}},
{{11'sd916, 8'sd-96, 12'sd1532}, {13'sd-2402, 13'sd2832, 13'sd-2789}, {12'sd1341, 12'sd1714, 13'sd-2761}},
{{12'sd1031, 12'sd1643, 12'sd-1304}, {11'sd653, 11'sd-867, 12'sd1437}, {12'sd-1221, 12'sd-1270, 12'sd1247}},
{{12'sd-2028, 11'sd-570, 12'sd1162}, {12'sd-1739, 11'sd-924, 12'sd1608}, {11'sd745, 11'sd1001, 12'sd-1158}}},
{
{{11'sd544, 12'sd1134, 12'sd1570}, {12'sd-1960, 12'sd1251, 11'sd718}, {9'sd143, 11'sd938, 12'sd1393}},
{{10'sd-397, 11'sd-745, 11'sd592}, {9'sd-223, 12'sd1986, 13'sd-2272}, {11'sd-918, 13'sd-3077, 12'sd1267}},
{{12'sd1187, 14'sd4393, 13'sd2807}, {13'sd2579, 13'sd3166, 13'sd2735}, {13'sd-2564, 11'sd-954, 13'sd-2944}},
{{11'sd755, 10'sd-439, 10'sd264}, {11'sd515, 12'sd-1056, 10'sd-368}, {10'sd-347, 10'sd345, 10'sd378}},
{{12'sd-1720, 8'sd-117, 12'sd-1801}, {12'sd1864, 13'sd-2141, 13'sd-2868}, {11'sd624, 11'sd-767, 12'sd-1924}},
{{11'sd703, 13'sd2660, 12'sd1658}, {13'sd-2523, 13'sd2134, 12'sd1753}, {13'sd2698, 12'sd-1588, 10'sd509}},
{{13'sd2473, 13'sd-2123, 11'sd1009}, {10'sd-428, 11'sd-835, 13'sd-2300}, {14'sd4756, 13'sd2845, 10'sd-313}},
{{12'sd1767, 11'sd862, 10'sd-411}, {11'sd785, 11'sd819, 12'sd-1872}, {8'sd-70, 12'sd1480, 13'sd-3160}},
{{13'sd3576, 11'sd612, 9'sd168}, {11'sd-731, 9'sd-156, 13'sd-3751}, {11'sd-556, 13'sd3287, 12'sd1204}},
{{13'sd2176, 13'sd2621, 9'sd-149}, {10'sd-358, 12'sd-1170, 11'sd-760}, {11'sd-876, 12'sd1716, 10'sd-295}},
{{12'sd-1769, 12'sd1961, 9'sd-229}, {7'sd-37, 10'sd-287, 13'sd-2238}, {12'sd-1305, 12'sd1958, 11'sd-594}},
{{12'sd1563, 8'sd70, 11'sd778}, {13'sd-3194, 13'sd-2127, 12'sd1273}, {12'sd-1325, 11'sd-854, 13'sd2687}},
{{12'sd2006, 13'sd-2690, 12'sd-1115}, {11'sd-838, 12'sd-1945, 12'sd1480}, {11'sd694, 12'sd1752, 12'sd-1110}},
{{12'sd-1242, 12'sd-1902, 12'sd-1103}, {12'sd1485, 12'sd1226, 10'sd320}, {12'sd1038, 13'sd2232, 13'sd2370}},
{{11'sd854, 13'sd2181, 11'sd783}, {10'sd-476, 10'sd-509, 13'sd-2126}, {13'sd-3263, 12'sd-1866, 13'sd-3474}},
{{13'sd-2736, 12'sd-1128, 11'sd-798}, {12'sd-2001, 10'sd-360, 12'sd-1708}, {8'sd80, 9'sd-174, 10'sd-268}},
{{10'sd300, 12'sd1440, 12'sd-1165}, {12'sd-1371, 13'sd2920, 12'sd1259}, {9'sd-228, 12'sd-1681, 10'sd-397}},
{{10'sd330, 11'sd-800, 13'sd-2263}, {12'sd-1195, 13'sd-2886, 9'sd-191}, {9'sd158, 13'sd-2807, 13'sd-3105}},
{{11'sd-851, 9'sd235, 9'sd183}, {12'sd1930, 10'sd280, 13'sd-2544}, {12'sd1803, 12'sd1549, 8'sd-68}},
{{11'sd-859, 11'sd-799, 11'sd-993}, {11'sd547, 13'sd-2194, 12'sd-1756}, {10'sd-445, 13'sd2818, 13'sd2749}},
{{12'sd1690, 13'sd2129, 13'sd3125}, {9'sd133, 13'sd-2541, 12'sd1347}, {13'sd3579, 7'sd-33, 12'sd1061}},
{{12'sd-1223, 13'sd-2170, 9'sd250}, {11'sd-1016, 9'sd190, 11'sd-733}, {11'sd-699, 12'sd1154, 9'sd-151}},
{{13'sd-2200, 11'sd-740, 13'sd2187}, {12'sd-1291, 13'sd-2555, 12'sd-1478}, {13'sd-2633, 12'sd-1336, 12'sd-1565}},
{{13'sd2513, 13'sd2262, 11'sd570}, {13'sd2241, 11'sd649, 12'sd-1329}, {13'sd2133, 12'sd-1316, 10'sd350}},
{{12'sd1530, 12'sd-1899, 12'sd-1477}, {10'sd405, 12'sd1167, 11'sd-531}, {11'sd947, 10'sd-310, 8'sd-64}},
{{12'sd-1879, 11'sd-971, 8'sd-105}, {6'sd28, 12'sd1300, 12'sd-1079}, {12'sd-1168, 12'sd1109, 12'sd-1539}},
{{13'sd2203, 10'sd-321, 13'sd2078}, {11'sd872, 12'sd1535, 12'sd1893}, {12'sd-1378, 13'sd2142, 10'sd304}},
{{11'sd-835, 12'sd1175, 10'sd-430}, {11'sd976, 13'sd2683, 12'sd-1739}, {9'sd-234, 13'sd2372, 6'sd-22}},
{{12'sd-1220, 10'sd284, 13'sd2555}, {12'sd-1777, 10'sd-481, 12'sd-1030}, {13'sd-2897, 7'sd61, 11'sd655}},
{{12'sd-1149, 12'sd-1505, 10'sd-339}, {13'sd2182, 13'sd-2763, 13'sd-2268}, {11'sd-859, 11'sd-533, 9'sd241}},
{{6'sd-22, 12'sd1794, 11'sd754}, {12'sd1544, 13'sd2129, 13'sd2448}, {11'sd800, 13'sd3575, 11'sd552}},
{{12'sd-1744, 13'sd2761, 13'sd2659}, {12'sd-1339, 10'sd-405, 12'sd-1895}, {11'sd821, 12'sd1477, 9'sd-197}},
{{13'sd-2707, 13'sd-3317, 13'sd-2306}, {10'sd-284, 10'sd386, 10'sd376}, {9'sd-195, 12'sd1383, 11'sd-823}},
{{13'sd2844, 13'sd2518, 12'sd-1624}, {13'sd3403, 12'sd1245, 11'sd-578}, {13'sd-2366, 13'sd-2662, 12'sd-1184}},
{{12'sd1307, 12'sd1818, 12'sd1857}, {13'sd2632, 12'sd1166, 13'sd3276}, {11'sd901, 13'sd2809, 11'sd678}},
{{8'sd79, 12'sd-1989, 11'sd-671}, {11'sd618, 11'sd732, 10'sd-435}, {12'sd-2021, 12'sd1759, 11'sd940}},
{{11'sd987, 12'sd1954, 12'sd-1694}, {12'sd1329, 9'sd197, 10'sd464}, {9'sd186, 13'sd2643, 5'sd-15}},
{{13'sd-2499, 13'sd-2290, 12'sd-1840}, {13'sd2547, 13'sd2107, 12'sd-1961}, {10'sd429, 13'sd2949, 12'sd-1650}},
{{10'sd-447, 12'sd-1598, 11'sd880}, {10'sd-304, 11'sd-570, 12'sd1847}, {12'sd-1192, 13'sd-2504, 13'sd-2245}},
{{11'sd-582, 11'sd-760, 12'sd-1210}, {11'sd603, 11'sd-540, 10'sd443}, {11'sd-930, 13'sd-3366, 12'sd1561}},
{{10'sd-304, 12'sd1397, 12'sd-1375}, {10'sd375, 12'sd1903, 14'sd-4169}, {12'sd1802, 10'sd259, 13'sd2619}},
{{11'sd990, 11'sd-787, 13'sd3493}, {11'sd-585, 11'sd577, 10'sd-493}, {13'sd-2379, 12'sd-1998, 12'sd-1834}},
{{12'sd1879, 12'sd1181, 11'sd958}, {10'sd-323, 13'sd2741, 3'sd3}, {11'sd682, 13'sd3840, 12'sd1767}},
{{13'sd2065, 13'sd2312, 12'sd1986}, {12'sd1465, 12'sd1263, 12'sd1237}, {8'sd110, 12'sd-1466, 11'sd819}},
{{12'sd1376, 10'sd-421, 13'sd-2571}, {12'sd1236, 9'sd-139, 12'sd-1207}, {12'sd-1221, 13'sd2778, 11'sd-572}},
{{10'sd-323, 11'sd-563, 12'sd1708}, {13'sd2050, 12'sd-1803, 12'sd-1186}, {12'sd-1962, 12'sd-1102, 13'sd-2239}},
{{13'sd-2481, 11'sd-575, 11'sd-639}, {12'sd-1032, 10'sd307, 10'sd317}, {12'sd1416, 12'sd1295, 12'sd1527}},
{{13'sd3699, 13'sd2073, 12'sd1414}, {13'sd3521, 12'sd-1594, 12'sd-1350}, {12'sd-1569, 13'sd2715, 9'sd142}},
{{13'sd2066, 12'sd1114, 13'sd-3259}, {13'sd3461, 11'sd-929, 13'sd-3096}, {12'sd1352, 12'sd-1159, 8'sd-90}},
{{13'sd-2309, 14'sd-4720, 14'sd-4766}, {12'sd-1804, 12'sd1762, 5'sd8}, {6'sd30, 13'sd-2840, 14'sd-4733}},
{{12'sd-1106, 13'sd2340, 12'sd-1551}, {13'sd-3821, 11'sd-840, 12'sd-1582}, {10'sd-290, 10'sd-379, 11'sd823}},
{{8'sd84, 13'sd-2306, 11'sd-698}, {8'sd70, 12'sd-1111, 13'sd2472}, {12'sd1834, 11'sd-687, 9'sd-197}},
{{11'sd739, 12'sd1722, 10'sd-449}, {13'sd-2861, 12'sd-1319, 12'sd-1856}, {9'sd-176, 13'sd2056, 13'sd-2212}},
{{12'sd-1837, 12'sd1206, 12'sd1832}, {12'sd1286, 12'sd-1123, 11'sd839}, {6'sd29, 13'sd2291, 12'sd1790}},
{{12'sd-1127, 12'sd1442, 10'sd-462}, {12'sd-1431, 12'sd-1142, 12'sd1241}, {9'sd196, 13'sd-3072, 11'sd-632}},
{{12'sd1148, 11'sd657, 12'sd1584}, {12'sd-1885, 12'sd1700, 9'sd242}, {11'sd729, 13'sd3182, 12'sd1709}},
{{12'sd-1117, 6'sd28, 13'sd2297}, {11'sd-635, 13'sd-2050, 10'sd-375}, {9'sd169, 13'sd-2167, 13'sd-3064}},
{{11'sd834, 12'sd1829, 9'sd173}, {13'sd3531, 10'sd-469, 12'sd1532}, {12'sd1456, 13'sd-2205, 13'sd-2518}},
{{12'sd-2001, 13'sd-2355, 12'sd-1700}, {12'sd1135, 13'sd-2258, 12'sd-1957}, {12'sd1490, 11'sd1013, 7'sd-32}},
{{14'sd4133, 11'sd692, 14'sd4645}, {11'sd-659, 13'sd3626, 13'sd3490}, {14'sd4124, 13'sd2983, 13'sd2696}},
{{11'sd-851, 12'sd1582, 13'sd-2661}, {12'sd1501, 12'sd-1547, 13'sd-2925}, {12'sd1793, 11'sd-623, 11'sd719}},
{{13'sd-2309, 10'sd389, 10'sd263}, {9'sd205, 12'sd-1566, 13'sd2634}, {9'sd-209, 13'sd-2894, 9'sd142}},
{{13'sd2660, 11'sd-804, 13'sd3228}, {12'sd1734, 13'sd-2390, 12'sd-1174}, {12'sd1943, 13'sd2539, 13'sd2306}},
{{11'sd607, 13'sd2725, 11'sd661}, {11'sd950, 12'sd1804, 13'sd-2235}, {11'sd-987, 11'sd-911, 13'sd-3202}}},
{
{{12'sd-1792, 9'sd252, 13'sd2145}, {12'sd-1621, 12'sd1854, 11'sd637}, {11'sd-761, 13'sd-2107, 9'sd196}},
{{8'sd-66, 13'sd2633, 12'sd1391}, {12'sd1441, 13'sd-2251, 8'sd-74}, {11'sd-592, 12'sd-1877, 12'sd-1098}},
{{12'sd1519, 12'sd1851, 12'sd1529}, {13'sd2331, 13'sd-2821, 12'sd-1610}, {11'sd-995, 12'sd1231, 12'sd1198}},
{{11'sd-609, 11'sd-959, 11'sd-700}, {12'sd-1911, 12'sd-1697, 13'sd2790}, {13'sd-2334, 12'sd1044, 12'sd1592}},
{{11'sd-782, 12'sd1535, 12'sd1810}, {9'sd152, 9'sd-225, 11'sd-704}, {13'sd2261, 13'sd-2368, 12'sd1258}},
{{12'sd-1947, 11'sd911, 8'sd69}, {12'sd-1411, 12'sd-2003, 12'sd1274}, {12'sd1398, 12'sd-1220, 12'sd1074}},
{{12'sd1572, 12'sd1456, 13'sd-2198}, {11'sd-822, 12'sd1615, 8'sd-114}, {10'sd-508, 12'sd1949, 12'sd1054}},
{{13'sd-2786, 12'sd1907, 11'sd-554}, {13'sd2320, 10'sd413, 10'sd-402}, {8'sd114, 9'sd140, 12'sd1572}},
{{10'sd-460, 13'sd-2360, 12'sd-1105}, {11'sd546, 13'sd2252, 12'sd-1629}, {12'sd-1317, 12'sd-1384, 12'sd1692}},
{{11'sd-971, 10'sd330, 9'sd-235}, {12'sd-1271, 11'sd-961, 13'sd2667}, {6'sd20, 13'sd2298, 12'sd-1082}},
{{12'sd1453, 12'sd2022, 10'sd478}, {11'sd-914, 12'sd1852, 12'sd-1759}, {12'sd1388, 11'sd806, 10'sd359}},
{{11'sd-734, 8'sd93, 11'sd-737}, {13'sd-2645, 13'sd2319, 13'sd-2415}, {11'sd-791, 13'sd-2792, 13'sd-2211}},
{{12'sd-2040, 10'sd-365, 11'sd-766}, {12'sd-1050, 12'sd1239, 12'sd-1987}, {12'sd-2038, 12'sd-1220, 13'sd-2435}},
{{11'sd712, 11'sd-1004, 13'sd-2231}, {12'sd-1720, 12'sd-1792, 12'sd-1877}, {12'sd1342, 11'sd-860, 11'sd601}},
{{12'sd-1372, 12'sd-1296, 12'sd-1208}, {12'sd-1381, 10'sd297, 10'sd-509}, {13'sd-2233, 10'sd-293, 12'sd-1904}},
{{10'sd292, 13'sd2999, 12'sd-1541}, {10'sd-340, 13'sd2107, 13'sd-2192}, {13'sd-2591, 12'sd1573, 12'sd-1456}},
{{12'sd-1693, 10'sd-485, 11'sd712}, {9'sd222, 13'sd-2761, 12'sd1726}, {12'sd-1277, 13'sd2708, 12'sd-1635}},
{{13'sd3379, 12'sd1962, 11'sd-806}, {11'sd-868, 13'sd2855, 11'sd-967}, {13'sd-2186, 12'sd1726, 13'sd-2257}},
{{11'sd-1017, 10'sd288, 12'sd-1095}, {12'sd1296, 7'sd-53, 12'sd-1872}, {12'sd-1784, 12'sd-1246, 12'sd1325}},
{{11'sd-843, 12'sd1094, 12'sd1798}, {12'sd-2020, 11'sd1008, 12'sd-1659}, {12'sd1417, 6'sd-25, 8'sd-65}},
{{11'sd600, 12'sd1445, 11'sd-942}, {13'sd2059, 13'sd-2655, 11'sd-821}, {12'sd-1322, 11'sd-525, 13'sd2738}},
{{12'sd1786, 13'sd2343, 11'sd820}, {12'sd1886, 12'sd1842, 12'sd-1137}, {13'sd-2825, 13'sd-2316, 12'sd-1641}},
{{13'sd-2417, 11'sd968, 12'sd1646}, {12'sd-2036, 13'sd2434, 11'sd-695}, {12'sd1158, 12'sd1754, 12'sd1470}},
{{10'sd508, 13'sd-2100, 13'sd-2628}, {11'sd700, 13'sd-2609, 12'sd-1403}, {12'sd-1136, 12'sd1949, 12'sd1282}},
{{13'sd2526, 11'sd-696, 13'sd2468}, {10'sd-381, 10'sd414, 12'sd-1991}, {11'sd-567, 12'sd1570, 12'sd-1586}},
{{13'sd-2304, 12'sd1403, 12'sd1680}, {10'sd282, 13'sd2678, 10'sd304}, {9'sd-185, 12'sd1692, 12'sd-1951}},
{{13'sd-2620, 13'sd2276, 12'sd-1890}, {12'sd-1740, 13'sd-2938, 7'sd56}, {13'sd-2710, 12'sd-1183, 12'sd-1467}},
{{5'sd-15, 12'sd-1380, 13'sd-2441}, {13'sd2736, 10'sd-305, 12'sd1075}, {12'sd-1192, 12'sd-1994, 11'sd617}},
{{13'sd2609, 11'sd806, 12'sd1598}, {12'sd1727, 12'sd-1905, 8'sd-64}, {13'sd2477, 13'sd2197, 8'sd123}},
{{11'sd-906, 12'sd-1142, 10'sd441}, {11'sd904, 12'sd1979, 12'sd2041}, {12'sd-1199, 9'sd156, 8'sd-105}},
{{12'sd1080, 13'sd2923, 12'sd1764}, {13'sd2169, 8'sd-72, 8'sd-72}, {8'sd-111, 12'sd-1651, 13'sd-2456}},
{{10'sd-400, 13'sd2094, 12'sd-1338}, {13'sd2587, 10'sd270, 13'sd2267}, {10'sd-464, 13'sd2129, 12'sd-1427}},
{{12'sd-1897, 12'sd1188, 13'sd-2292}, {13'sd2648, 13'sd-2957, 11'sd-570}, {11'sd-734, 13'sd2216, 13'sd2395}},
{{10'sd440, 13'sd-2180, 13'sd2276}, {12'sd-1344, 8'sd-71, 13'sd2529}, {12'sd1096, 12'sd1775, 12'sd-1440}},
{{12'sd1967, 8'sd123, 11'sd-859}, {12'sd-1933, 10'sd-308, 12'sd-1458}, {9'sd157, 9'sd192, 13'sd-2648}},
{{13'sd-2092, 11'sd-575, 11'sd-643}, {12'sd1220, 11'sd656, 12'sd1716}, {12'sd1749, 12'sd1220, 12'sd2005}},
{{11'sd-950, 11'sd954, 13'sd2502}, {13'sd2134, 11'sd715, 13'sd2331}, {13'sd-2441, 12'sd1996, 13'sd2846}},
{{12'sd1889, 6'sd17, 13'sd-2283}, {12'sd1333, 13'sd2093, 11'sd-542}, {11'sd-670, 13'sd2484, 12'sd-1976}},
{{11'sd-514, 12'sd1664, 12'sd1900}, {11'sd819, 8'sd83, 12'sd-1367}, {13'sd2206, 13'sd-2591, 12'sd1489}},
{{12'sd1686, 11'sd982, 13'sd2539}, {11'sd-715, 12'sd-1805, 10'sd-331}, {11'sd-715, 12'sd1977, 13'sd2926}},
{{12'sd-1863, 12'sd-1800, 13'sd-3520}, {13'sd-3020, 11'sd969, 13'sd-2551}, {11'sd805, 11'sd715, 8'sd-96}},
{{12'sd-1581, 11'sd-927, 10'sd296}, {12'sd2009, 11'sd828, 13'sd-2052}, {13'sd-2557, 11'sd579, 6'sd23}},
{{12'sd-1927, 13'sd-2603, 12'sd1130}, {13'sd-2166, 11'sd-768, 12'sd-1033}, {13'sd-2844, 13'sd2131, 12'sd1918}},
{{10'sd290, 12'sd1182, 7'sd57}, {13'sd2232, 9'sd237, 11'sd920}, {11'sd980, 11'sd-1010, 11'sd-907}},
{{12'sd1500, 10'sd372, 12'sd1894}, {8'sd101, 11'sd-834, 13'sd2205}, {10'sd-392, 13'sd-2932, 13'sd2127}},
{{12'sd-1923, 10'sd-299, 11'sd797}, {12'sd-1665, 12'sd-1950, 13'sd3025}, {11'sd766, 12'sd-1197, 13'sd2703}},
{{13'sd2145, 13'sd-2059, 13'sd-2243}, {10'sd417, 13'sd2230, 12'sd1028}, {13'sd-2203, 13'sd-2354, 11'sd854}},
{{12'sd1686, 13'sd2614, 11'sd728}, {13'sd-2575, 11'sd835, 12'sd1895}, {13'sd-3087, 12'sd1624, 10'sd272}},
{{11'sd-1021, 13'sd-2095, 13'sd2502}, {11'sd-793, 12'sd1878, 9'sd179}, {10'sd379, 13'sd3710, 11'sd860}},
{{13'sd-2459, 12'sd1484, 13'sd-2660}, {10'sd-363, 10'sd-277, 8'sd-74}, {12'sd1279, 13'sd3484, 12'sd-1559}},
{{11'sd587, 11'sd788, 12'sd-1839}, {8'sd-95, 13'sd-2317, 11'sd914}, {13'sd2554, 10'sd-436, 12'sd-1462}},
{{11'sd-687, 12'sd2003, 12'sd-1033}, {13'sd2706, 9'sd-180, 12'sd-1174}, {12'sd1036, 11'sd976, 11'sd-996}},
{{11'sd-557, 13'sd2524, 13'sd2534}, {13'sd-2537, 11'sd-872, 12'sd-1089}, {11'sd764, 11'sd-759, 10'sd399}},
{{12'sd1707, 13'sd-2840, 8'sd75}, {13'sd2142, 13'sd-2994, 11'sd562}, {9'sd145, 12'sd-1357, 13'sd-2537}},
{{13'sd2633, 12'sd1777, 10'sd-410}, {12'sd-1233, 10'sd323, 12'sd-1185}, {11'sd-583, 7'sd54, 11'sd533}},
{{11'sd-587, 12'sd1905, 13'sd-2497}, {12'sd1812, 12'sd1408, 11'sd900}, {12'sd-1730, 13'sd-2050, 11'sd-740}},
{{9'sd-233, 12'sd1935, 10'sd-274}, {8'sd-81, 12'sd1660, 12'sd-1541}, {10'sd-414, 10'sd-469, 13'sd2468}},
{{12'sd-1716, 8'sd76, 9'sd141}, {10'sd401, 12'sd-1947, 9'sd-178}, {12'sd-1747, 11'sd862, 8'sd-79}},
{{12'sd-1858, 11'sd-930, 12'sd-1985}, {13'sd-2076, 11'sd575, 11'sd568}, {12'sd-1163, 12'sd1220, 11'sd-812}},
{{13'sd2975, 13'sd2573, 12'sd1152}, {13'sd-2709, 10'sd502, 11'sd-976}, {13'sd-2988, 13'sd-2478, 10'sd-438}},
{{12'sd-1581, 12'sd-1817, 10'sd-425}, {13'sd2347, 1'sd0, 13'sd2095}, {11'sd-642, 13'sd2468, 11'sd1012}},
{{12'sd1997, 13'sd2573, 13'sd-2449}, {8'sd-115, 9'sd-136, 13'sd-2190}, {13'sd2461, 12'sd-1569, 11'sd966}},
{{13'sd3343, 10'sd-460, 12'sd2022}, {12'sd-1324, 13'sd-2097, 8'sd-114}, {10'sd-367, 5'sd-9, 13'sd-2282}},
{{12'sd1305, 12'sd1212, 8'sd121}, {12'sd1234, 11'sd1011, 13'sd2240}, {13'sd-2066, 12'sd-1403, 10'sd-421}}},
{
{{12'sd1452, 13'sd-2269, 12'sd1138}, {11'sd-972, 12'sd-1529, 11'sd688}, {12'sd1942, 13'sd-2283, 13'sd-2112}},
{{11'sd972, 8'sd-122, 12'sd2002}, {12'sd1272, 12'sd-1407, 13'sd-2245}, {12'sd1680, 10'sd358, 12'sd-1641}},
{{13'sd-3787, 12'sd-1450, 11'sd958}, {12'sd1162, 11'sd-624, 11'sd513}, {13'sd-3771, 10'sd-261, 13'sd-3237}},
{{11'sd875, 11'sd516, 11'sd-525}, {9'sd-156, 12'sd1542, 12'sd1035}, {13'sd2557, 13'sd-2246, 11'sd-883}},
{{11'sd-560, 13'sd-2814, 13'sd2053}, {11'sd872, 12'sd1740, 10'sd406}, {6'sd-23, 9'sd228, 12'sd1247}},
{{12'sd-1692, 13'sd-2181, 10'sd473}, {9'sd146, 11'sd-865, 12'sd1056}, {12'sd1314, 13'sd2172, 12'sd1108}},
{{11'sd-788, 12'sd-1264, 13'sd-2090}, {12'sd1641, 12'sd1174, 12'sd-1090}, {9'sd206, 12'sd-1108, 13'sd3391}},
{{12'sd1577, 12'sd-1741, 13'sd-3432}, {13'sd2913, 12'sd1161, 8'sd113}, {12'sd-1954, 11'sd556, 11'sd677}},
{{10'sd-367, 12'sd1439, 12'sd-1821}, {12'sd-1674, 13'sd-2573, 13'sd-3275}, {11'sd-744, 13'sd-2830, 12'sd1933}},
{{12'sd1414, 11'sd653, 13'sd-2538}, {13'sd2209, 12'sd-1321, 12'sd-1889}, {13'sd2865, 12'sd1071, 13'sd-2419}},
{{13'sd-2077, 13'sd-2370, 9'sd-212}, {10'sd312, 11'sd528, 11'sd-927}, {12'sd1151, 13'sd-2130, 11'sd-969}},
{{12'sd-1643, 13'sd2846, 11'sd-756}, {11'sd-801, 11'sd-602, 12'sd1429}, {13'sd2603, 11'sd594, 11'sd541}},
{{11'sd913, 13'sd2145, 10'sd-438}, {11'sd739, 12'sd-1382, 7'sd-40}, {13'sd3488, 13'sd3657, 13'sd3444}},
{{10'sd-265, 12'sd1547, 12'sd-1702}, {12'sd-1139, 11'sd782, 12'sd-1677}, {13'sd-2094, 9'sd-192, 12'sd-1980}},
{{11'sd725, 10'sd-450, 12'sd-1105}, {13'sd2169, 12'sd1884, 13'sd-2345}, {12'sd-1807, 10'sd336, 13'sd-2728}},
{{11'sd544, 12'sd1071, 12'sd-2010}, {8'sd124, 13'sd-2406, 12'sd-1743}, {10'sd-295, 12'sd-2021, 12'sd-1137}},
{{11'sd700, 13'sd2458, 12'sd1711}, {12'sd-1376, 12'sd-1278, 12'sd-1515}, {12'sd1913, 12'sd-1831, 12'sd-1697}},
{{10'sd-334, 12'sd1630, 12'sd1541}, {13'sd2438, 11'sd936, 13'sd2263}, {8'sd89, 11'sd540, 13'sd2584}},
{{10'sd316, 12'sd1036, 10'sd385}, {8'sd-82, 11'sd-873, 12'sd1753}, {12'sd-1070, 12'sd-1550, 13'sd-2528}},
{{13'sd-2140, 10'sd-415, 13'sd-2243}, {9'sd-248, 13'sd-2241, 13'sd-2589}, {11'sd-916, 11'sd799, 12'sd1396}},
{{7'sd-56, 7'sd-56, 12'sd1893}, {12'sd-1525, 10'sd-275, 13'sd2556}, {12'sd1268, 11'sd583, 12'sd-1049}},
{{12'sd-1330, 13'sd-3013, 12'sd1113}, {12'sd1930, 12'sd1177, 13'sd2052}, {12'sd-1242, 9'sd232, 12'sd1287}},
{{13'sd-2409, 13'sd2205, 11'sd-733}, {13'sd2233, 12'sd1409, 11'sd-934}, {12'sd1439, 13'sd-2656, 12'sd1207}},
{{11'sd650, 13'sd2566, 12'sd-1068}, {13'sd2780, 11'sd-551, 11'sd-581}, {13'sd2146, 12'sd1625, 12'sd-1972}},
{{10'sd-406, 12'sd-1550, 10'sd-344}, {13'sd2544, 12'sd-1287, 13'sd2272}, {12'sd1763, 13'sd2251, 11'sd-723}},
{{13'sd-2787, 11'sd751, 12'sd1863}, {12'sd-1263, 8'sd-121, 11'sd649}, {12'sd1183, 6'sd29, 11'sd779}},
{{12'sd1590, 11'sd-740, 11'sd851}, {13'sd-2111, 13'sd-2381, 13'sd-2467}, {12'sd-1351, 11'sd-974, 13'sd-2284}},
{{9'sd245, 13'sd-2840, 12'sd-1744}, {11'sd-978, 5'sd9, 12'sd-1633}, {10'sd478, 11'sd-817, 12'sd1042}},
{{12'sd1340, 12'sd1358, 11'sd844}, {12'sd1613, 13'sd2172, 12'sd1061}, {13'sd-2654, 13'sd2382, 10'sd-369}},
{{13'sd2263, 7'sd-57, 11'sd-997}, {13'sd2666, 13'sd2316, 13'sd-2216}, {12'sd1190, 13'sd2579, 12'sd1590}},
{{10'sd256, 13'sd2404, 10'sd382}, {13'sd2383, 11'sd-533, 9'sd-209}, {12'sd1250, 14'sd4386, 9'sd135}},
{{12'sd-1323, 12'sd-1849, 13'sd2382}, {12'sd1488, 12'sd-1372, 12'sd1031}, {11'sd-550, 12'sd1074, 13'sd2057}},
{{13'sd3118, 13'sd2563, 11'sd-591}, {13'sd2328, 11'sd764, 11'sd834}, {14'sd4176, 12'sd-1299, 9'sd-250}},
{{13'sd-2597, 10'sd338, 9'sd-235}, {11'sd773, 13'sd2960, 12'sd1457}, {13'sd-3613, 12'sd1238, 12'sd-1629}},
{{12'sd-1189, 12'sd-1421, 13'sd-2266}, {12'sd1925, 11'sd528, 13'sd2475}, {12'sd-1484, 11'sd-656, 12'sd1904}},
{{13'sd2374, 12'sd1507, 13'sd2106}, {13'sd2287, 12'sd-1982, 8'sd65}, {9'sd-250, 9'sd131, 13'sd2638}},
{{11'sd765, 7'sd-61, 12'sd-1736}, {13'sd2654, 13'sd-2340, 13'sd2247}, {12'sd1695, 12'sd-1214, 11'sd-775}},
{{9'sd252, 13'sd-2316, 12'sd1780}, {13'sd2344, 10'sd459, 13'sd2804}, {12'sd1182, 7'sd37, 11'sd674}},
{{12'sd1233, 10'sd-368, 12'sd1157}, {10'sd-328, 13'sd2335, 12'sd1422}, {10'sd-295, 13'sd3292, 12'sd1337}},
{{12'sd1243, 12'sd1367, 12'sd-1466}, {12'sd1508, 13'sd2721, 8'sd-91}, {13'sd2975, 12'sd1617, 10'sd265}},
{{12'sd-1132, 12'sd1626, 11'sd-878}, {12'sd1032, 13'sd2202, 12'sd1340}, {10'sd-326, 11'sd810, 10'sd429}},
{{9'sd208, 13'sd-3482, 13'sd-2253}, {12'sd-1961, 10'sd274, 12'sd-1780}, {11'sd-688, 10'sd461, 12'sd1278}},
{{12'sd1782, 11'sd954, 13'sd2561}, {12'sd1176, 13'sd-2781, 11'sd594}, {12'sd-1630, 9'sd-162, 11'sd-797}},
{{13'sd2376, 13'sd-2204, 13'sd2275}, {12'sd1841, 12'sd1488, 11'sd-706}, {12'sd1461, 12'sd1838, 10'sd-385}},
{{12'sd-1754, 13'sd-2205, 9'sd213}, {12'sd1857, 12'sd-1612, 12'sd1479}, {12'sd-1952, 12'sd1592, 11'sd-566}},
{{5'sd-11, 11'sd677, 12'sd1335}, {9'sd-207, 11'sd-615, 12'sd1638}, {11'sd817, 13'sd-2219, 13'sd-2232}},
{{8'sd68, 12'sd1686, 12'sd1193}, {13'sd-2102, 11'sd767, 13'sd-2301}, {13'sd2108, 11'sd-650, 6'sd-17}},
{{13'sd-3087, 10'sd-460, 11'sd570}, {12'sd1433, 13'sd2783, 13'sd2773}, {12'sd2033, 7'sd-43, 11'sd-860}},
{{13'sd3247, 8'sd75, 11'sd909}, {13'sd2851, 13'sd-2905, 10'sd-411}, {7'sd61, 12'sd-1569, 11'sd-918}},
{{10'sd322, 8'sd-64, 10'sd-502}, {13'sd-3163, 13'sd-2756, 13'sd-2114}, {13'sd2569, 8'sd-75, 12'sd1132}},
{{12'sd-1976, 11'sd609, 13'sd2142}, {9'sd134, 11'sd-930, 13'sd2074}, {13'sd2987, 11'sd844, 13'sd2462}},
{{13'sd-2162, 12'sd1066, 13'sd2308}, {11'sd554, 13'sd-2201, 13'sd-2281}, {11'sd-969, 12'sd-1844, 11'sd-658}},
{{12'sd-1857, 12'sd-1134, 11'sd829}, {12'sd-1842, 12'sd-1600, 12'sd1756}, {11'sd855, 12'sd1979, 10'sd476}},
{{12'sd-1139, 13'sd-2736, 13'sd2274}, {12'sd-2000, 9'sd187, 12'sd-1201}, {13'sd-2387, 13'sd2326, 12'sd1403}},
{{12'sd-1085, 8'sd-98, 13'sd-4025}, {13'sd2192, 13'sd2171, 13'sd3250}, {11'sd731, 12'sd-1189, 12'sd-1210}},
{{12'sd1767, 13'sd-2250, 12'sd1105}, {10'sd-331, 12'sd-1444, 12'sd-1111}, {13'sd2352, 12'sd-1976, 11'sd-1008}},
{{12'sd-1233, 12'sd1927, 12'sd1969}, {10'sd-462, 9'sd-224, 10'sd292}, {12'sd1252, 11'sd-570, 12'sd1456}},
{{13'sd-3315, 13'sd-2114, 13'sd-3762}, {12'sd-1992, 13'sd2107, 12'sd-1872}, {14'sd-4512, 13'sd-3513, 12'sd-1934}},
{{10'sd-314, 12'sd1404, 13'sd2463}, {9'sd-173, 12'sd1972, 13'sd2689}, {12'sd-1841, 12'sd1525, 12'sd-1083}},
{{9'sd-246, 13'sd2476, 11'sd-898}, {10'sd440, 11'sd-967, 13'sd2854}, {12'sd-1519, 9'sd135, 11'sd787}},
{{13'sd-2584, 12'sd1189, 11'sd-649}, {13'sd-2362, 10'sd-430, 13'sd2401}, {12'sd1675, 9'sd245, 10'sd-448}},
{{12'sd-1700, 4'sd-4, 12'sd-1256}, {8'sd-111, 12'sd-1819, 11'sd-637}, {12'sd-1237, 10'sd-495, 12'sd1501}},
{{13'sd2617, 12'sd-1654, 13'sd-2185}, {12'sd-1553, 13'sd2957, 11'sd849}, {13'sd2202, 13'sd2401, 12'sd1820}},
{{11'sd1013, 12'sd1771, 13'sd-2218}, {11'sd858, 8'sd-69, 12'sd1572}, {13'sd2073, 11'sd864, 9'sd166}}},
{
{{10'sd-483, 12'sd1184, 11'sd-958}, {12'sd1362, 12'sd1567, 10'sd271}, {13'sd-3321, 10'sd-376, 12'sd-1962}},
{{13'sd-2903, 13'sd-2770, 13'sd-2412}, {13'sd-2618, 10'sd420, 11'sd-925}, {7'sd-62, 12'sd1477, 12'sd1931}},
{{12'sd-1441, 12'sd1515, 13'sd-2119}, {10'sd355, 11'sd657, 12'sd1821}, {12'sd-1501, 13'sd3769, 10'sd-331}},
{{7'sd46, 13'sd3076, 9'sd169}, {12'sd-1991, 11'sd849, 13'sd-2687}, {11'sd630, 9'sd-145, 13'sd-2332}},
{{10'sd303, 12'sd1268, 12'sd-1502}, {6'sd-31, 12'sd1186, 12'sd-1446}, {11'sd579, 10'sd-417, 12'sd-1118}},
{{9'sd191, 10'sd-318, 8'sd121}, {13'sd-2463, 13'sd2428, 8'sd-124}, {13'sd-2115, 3'sd-2, 12'sd1646}},
{{9'sd244, 10'sd-501, 12'sd2004}, {12'sd-1344, 12'sd-1409, 12'sd1287}, {12'sd1130, 12'sd1317, 11'sd918}},
{{9'sd156, 13'sd-2188, 10'sd268}, {13'sd2712, 12'sd-1571, 12'sd1215}, {13'sd-2052, 10'sd-288, 8'sd91}},
{{12'sd1647, 13'sd-2107, 11'sd-513}, {11'sd-797, 12'sd-1946, 8'sd111}, {9'sd-215, 12'sd1341, 13'sd-3085}},
{{13'sd2114, 12'sd-1366, 10'sd484}, {13'sd2150, 12'sd-1941, 11'sd-585}, {11'sd-553, 12'sd-1828, 9'sd245}},
{{12'sd-1616, 13'sd-2168, 12'sd1790}, {12'sd-1029, 12'sd1024, 13'sd-2647}, {13'sd2603, 12'sd1373, 13'sd-2171}},
{{13'sd-3064, 11'sd-773, 9'sd-180}, {12'sd-1726, 9'sd142, 13'sd2612}, {10'sd-468, 10'sd-387, 9'sd181}},
{{14'sd-6231, 11'sd538, 13'sd-2647}, {11'sd840, 11'sd-608, 13'sd3083}, {9'sd243, 13'sd2335, 13'sd3345}},
{{12'sd-1270, 11'sd768, 11'sd932}, {11'sd-561, 11'sd-710, 7'sd-51}, {11'sd-918, 12'sd-1545, 12'sd-1889}},
{{12'sd-1655, 11'sd-779, 11'sd-642}, {10'sd331, 12'sd1804, 13'sd-2426}, {12'sd-1965, 7'sd39, 12'sd-1517}},
{{10'sd-434, 7'sd-39, 11'sd850}, {12'sd-1895, 12'sd1078, 13'sd-2362}, {10'sd372, 12'sd-1156, 12'sd1235}},
{{11'sd711, 12'sd1430, 12'sd-1801}, {11'sd-957, 10'sd366, 13'sd-2610}, {13'sd-2291, 13'sd-2564, 13'sd-2905}},
{{10'sd-471, 13'sd-2666, 12'sd-1138}, {13'sd2876, 12'sd1358, 14'sd-4689}, {14'sd6075, 10'sd-318, 10'sd311}},
{{9'sd-232, 11'sd-951, 12'sd-1809}, {12'sd-1875, 11'sd874, 13'sd2075}, {12'sd1563, 13'sd3046, 10'sd-302}},
{{10'sd-467, 10'sd472, 12'sd-1321}, {9'sd-133, 12'sd1052, 12'sd-1333}, {12'sd1346, 13'sd-2242, 13'sd-2179}},
{{11'sd-948, 11'sd995, 12'sd-1192}, {13'sd2467, 11'sd660, 12'sd-1239}, {9'sd-236, 12'sd-1306, 13'sd-2988}},
{{12'sd-1851, 9'sd-194, 7'sd55}, {12'sd1440, 13'sd2770, 11'sd670}, {13'sd2546, 13'sd2198, 11'sd1000}},
{{11'sd876, 13'sd-2463, 12'sd-1456}, {11'sd-1003, 13'sd2657, 12'sd-1351}, {13'sd-2148, 8'sd95, 12'sd-1967}},
{{11'sd-878, 13'sd2139, 11'sd1013}, {9'sd-173, 12'sd-1208, 11'sd700}, {12'sd1905, 13'sd-2548, 11'sd-663}},
{{12'sd1702, 13'sd2990, 11'sd-741}, {12'sd-1385, 9'sd-152, 9'sd169}, {10'sd382, 12'sd-1086, 12'sd1166}},
{{5'sd-14, 11'sd-750, 11'sd565}, {13'sd-2069, 13'sd-2160, 10'sd-418}, {13'sd-2406, 12'sd-1369, 13'sd2203}},
{{10'sd-397, 13'sd2291, 13'sd2522}, {13'sd2891, 8'sd92, 11'sd-567}, {11'sd-600, 12'sd-1697, 11'sd563}},
{{11'sd-544, 13'sd-2854, 12'sd1202}, {12'sd1328, 12'sd1791, 12'sd-1280}, {11'sd632, 13'sd-3453, 12'sd-1654}},
{{12'sd-1236, 11'sd1005, 11'sd-778}, {11'sd816, 12'sd1463, 13'sd2547}, {13'sd2262, 10'sd-429, 13'sd2377}},
{{12'sd-1747, 11'sd-741, 9'sd229}, {13'sd-2089, 13'sd-2686, 9'sd188}, {13'sd2374, 12'sd1787, 12'sd1315}},
{{14'sd5417, 8'sd114, 12'sd-1659}, {14'sd5403, 12'sd-1070, 12'sd2005}, {14'sd6621, 9'sd-151, 12'sd1883}},
{{11'sd-558, 11'sd-660, 13'sd-3575}, {12'sd-1113, 10'sd373, 12'sd-1238}, {13'sd-2530, 13'sd-2410, 12'sd1701}},
{{13'sd2642, 12'sd-1146, 11'sd-1012}, {6'sd30, 12'sd-1740, 7'sd32}, {12'sd1816, 4'sd-4, 13'sd-2751}},
{{13'sd2981, 12'sd1608, 9'sd-169}, {13'sd2534, 13'sd-2656, 8'sd105}, {12'sd1724, 12'sd-1565, 12'sd1634}},
{{12'sd1153, 12'sd1811, 12'sd1451}, {8'sd87, 9'sd218, 12'sd1359}, {10'sd315, 11'sd-749, 11'sd-694}},
{{13'sd-2155, 12'sd1448, 9'sd-247}, {13'sd2295, 13'sd-2079, 12'sd-1384}, {12'sd-1519, 13'sd2510, 11'sd-542}},
{{12'sd-1947, 10'sd300, 12'sd-1263}, {11'sd-789, 13'sd-2153, 13'sd2117}, {12'sd1701, 12'sd1216, 12'sd1070}},
{{13'sd2397, 10'sd-449, 11'sd867}, {13'sd-2564, 13'sd-2241, 13'sd2644}, {12'sd1752, 9'sd202, 12'sd-1847}},
{{13'sd-3407, 5'sd14, 11'sd966}, {10'sd-458, 10'sd-471, 13'sd2705}, {12'sd1984, 13'sd-2438, 11'sd940}},
{{10'sd504, 12'sd1755, 9'sd198}, {10'sd417, 12'sd1058, 11'sd972}, {13'sd2462, 12'sd-1495, 12'sd1461}},
{{12'sd-1778, 12'sd1490, 11'sd651}, {13'sd-2621, 12'sd1123, 11'sd534}, {14'sd-4916, 12'sd-1709, 10'sd399}},
{{13'sd-3163, 11'sd-616, 7'sd-44}, {9'sd-221, 11'sd-1014, 10'sd-305}, {10'sd-393, 10'sd498, 9'sd194}},
{{12'sd1309, 13'sd2380, 13'sd2568}, {13'sd-3344, 11'sd534, 12'sd1132}, {13'sd-4068, 10'sd-359, 12'sd-1267}},
{{12'sd-1676, 8'sd119, 8'sd83}, {12'sd1363, 11'sd-891, 13'sd2468}, {13'sd-2456, 13'sd2301, 13'sd2401}},
{{12'sd-1990, 12'sd-1636, 13'sd2311}, {11'sd-646, 13'sd-2381, 12'sd-2042}, {13'sd-3398, 12'sd1825, 12'sd1948}},
{{11'sd883, 10'sd-349, 7'sd55}, {10'sd380, 13'sd-2233, 9'sd-181}, {11'sd544, 12'sd-1420, 11'sd-882}},
{{9'sd-173, 11'sd-598, 12'sd-1064}, {9'sd-186, 13'sd2479, 12'sd-1399}, {13'sd-2108, 8'sd102, 9'sd-131}},
{{12'sd-1206, 8'sd-122, 13'sd2370}, {13'sd2151, 13'sd3412, 13'sd2143}, {13'sd2176, 12'sd-1856, 13'sd3147}},
{{12'sd1640, 9'sd182, 12'sd1598}, {9'sd252, 9'sd-143, 13'sd-2900}, {13'sd2525, 13'sd-2530, 12'sd-1865}},
{{11'sd-786, 10'sd-504, 12'sd-1557}, {12'sd1105, 12'sd1786, 13'sd-2249}, {12'sd-1823, 11'sd786, 6'sd29}},
{{12'sd-1906, 13'sd2257, 11'sd-743}, {13'sd-2149, 13'sd-2363, 12'sd2036}, {13'sd-3249, 13'sd-2480, 12'sd1875}},
{{13'sd2287, 12'sd1308, 12'sd-1993}, {12'sd1335, 13'sd-2446, 11'sd-973}, {13'sd-2238, 8'sd89, 13'sd-2406}},
{{13'sd2366, 12'sd1161, 12'sd1386}, {10'sd509, 13'sd2277, 11'sd-612}, {13'sd2560, 11'sd736, 12'sd1240}},
{{8'sd-89, 12'sd1547, 12'sd1132}, {10'sd426, 12'sd1425, 12'sd-1994}, {9'sd188, 12'sd1394, 12'sd1896}},
{{10'sd-434, 13'sd-3777, 13'sd-2954}, {11'sd-832, 12'sd-1444, 12'sd-1405}, {13'sd2206, 11'sd-737, 12'sd1527}},
{{13'sd-2824, 9'sd143, 13'sd2281}, {10'sd-320, 11'sd703, 12'sd-1431}, {12'sd-1966, 12'sd1262, 13'sd2831}},
{{9'sd135, 12'sd1136, 12'sd1771}, {12'sd1922, 9'sd245, 12'sd-1889}, {12'sd1928, 11'sd822, 12'sd1871}},
{{5'sd15, 13'sd2476, 13'sd2653}, {12'sd-1980, 12'sd-1187, 13'sd2231}, {13'sd2824, 12'sd1873, 11'sd549}},
{{11'sd714, 12'sd-1967, 12'sd-1825}, {13'sd-2116, 12'sd1722, 10'sd-321}, {13'sd2622, 12'sd1429, 13'sd-2124}},
{{7'sd-63, 13'sd-2234, 9'sd-255}, {13'sd-2367, 12'sd-1268, 12'sd1156}, {11'sd810, 13'sd2172, 12'sd1857}},
{{10'sd308, 11'sd-923, 13'sd-2613}, {12'sd-1550, 12'sd-1896, 12'sd1493}, {12'sd1249, 8'sd122, 12'sd1978}},
{{12'sd1307, 11'sd958, 12'sd1902}, {13'sd2743, 11'sd-1015, 12'sd1760}, {13'sd2668, 12'sd-1889, 8'sd105}},
{{12'sd1860, 11'sd525, 13'sd2423}, {12'sd-1178, 13'sd2645, 13'sd3251}, {12'sd1430, 13'sd2950, 10'sd-371}},
{{12'sd1653, 13'sd-2928, 13'sd-2347}, {13'sd2907, 12'sd-1029, 11'sd-613}, {13'sd2944, 12'sd1277, 11'sd973}}},
{
{{11'sd-740, 10'sd486, 10'sd284}, {9'sd218, 13'sd-2536, 12'sd-1272}, {12'sd1146, 10'sd-288, 13'sd2322}},
{{13'sd3111, 12'sd-1438, 11'sd-719}, {12'sd1147, 13'sd-2535, 11'sd-724}, {13'sd2649, 11'sd-621, 12'sd1841}},
{{11'sd867, 10'sd491, 14'sd5437}, {13'sd-3357, 12'sd1677, 13'sd2561}, {12'sd-1063, 10'sd-408, 11'sd735}},
{{9'sd-212, 12'sd-1132, 12'sd1036}, {12'sd1367, 10'sd-395, 12'sd-1485}, {12'sd-1617, 11'sd606, 12'sd-1064}},
{{11'sd769, 11'sd964, 11'sd-911}, {13'sd2873, 13'sd2449, 12'sd-1678}, {13'sd2172, 12'sd-1393, 10'sd-453}},
{{12'sd1293, 11'sd-752, 11'sd693}, {12'sd1850, 9'sd214, 12'sd-1834}, {12'sd1970, 11'sd-837, 13'sd2716}},
{{9'sd132, 13'sd-2501, 11'sd542}, {11'sd843, 12'sd-1330, 11'sd-707}, {14'sd4153, 10'sd346, 12'sd1471}},
{{12'sd1529, 11'sd849, 13'sd2375}, {13'sd-2834, 12'sd1920, 13'sd2397}, {12'sd-1855, 12'sd-1878, 13'sd2078}},
{{10'sd284, 12'sd1677, 13'sd-3105}, {9'sd-133, 11'sd-674, 14'sd-4646}, {10'sd329, 12'sd-1066, 12'sd-1241}},
{{11'sd-725, 11'sd-1015, 12'sd2042}, {13'sd-2060, 12'sd-1122, 11'sd-1010}, {10'sd456, 13'sd2090, 11'sd787}},
{{12'sd-1972, 13'sd-2610, 11'sd-704}, {12'sd1210, 13'sd2492, 13'sd3237}, {12'sd-1821, 13'sd2136, 13'sd2623}},
{{13'sd2376, 9'sd184, 12'sd1660}, {13'sd-2495, 13'sd-2155, 12'sd-1611}, {13'sd-2173, 13'sd-2722, 13'sd-2117}},
{{10'sd477, 13'sd-2511, 11'sd844}, {12'sd1743, 13'sd-2407, 13'sd-2613}, {13'sd-3076, 13'sd-3946, 13'sd-3886}},
{{11'sd-948, 13'sd2648, 9'sd222}, {13'sd-2131, 9'sd-255, 12'sd-1738}, {11'sd725, 9'sd236, 13'sd-3016}},
{{11'sd-727, 12'sd-1775, 12'sd-1783}, {9'sd212, 13'sd-2369, 13'sd-3673}, {13'sd-2555, 13'sd2619, 11'sd607}},
{{13'sd-2203, 13'sd2819, 12'sd1498}, {13'sd-2285, 12'sd1520, 11'sd816}, {13'sd-3621, 12'sd-1862, 10'sd-498}},
{{10'sd-420, 12'sd1944, 10'sd287}, {13'sd2829, 13'sd3037, 13'sd2785}, {12'sd1447, 12'sd1820, 13'sd-2300}},
{{11'sd-858, 12'sd-1510, 12'sd1122}, {13'sd2697, 13'sd2986, 9'sd182}, {13'sd-2124, 13'sd-3469, 12'sd1056}},
{{12'sd1196, 13'sd-2468, 13'sd-2383}, {10'sd-283, 11'sd-725, 12'sd-1036}, {9'sd-228, 10'sd-488, 13'sd-2231}},
{{13'sd-2653, 13'sd-2331, 11'sd-570}, {13'sd-2427, 12'sd1719, 12'sd1610}, {11'sd-626, 12'sd-1309, 5'sd11}},
{{12'sd1422, 13'sd-2631, 13'sd2935}, {12'sd-1418, 13'sd2095, 12'sd1582}, {12'sd1927, 12'sd-1779, 13'sd2888}},
{{12'sd-1777, 11'sd-853, 12'sd1644}, {9'sd202, 12'sd1564, 11'sd951}, {11'sd758, 8'sd-89, 11'sd903}},
{{9'sd-245, 12'sd1837, 11'sd797}, {13'sd-2947, 12'sd-1746, 10'sd-372}, {13'sd-2955, 12'sd1969, 11'sd-654}},
{{12'sd1815, 8'sd73, 12'sd-1142}, {12'sd-2021, 12'sd1967, 11'sd645}, {11'sd-963, 12'sd1655, 13'sd2173}},
{{10'sd-364, 12'sd-1846, 7'sd-36}, {10'sd-308, 13'sd2172, 13'sd2886}, {12'sd-1783, 11'sd-767, 13'sd3004}},
{{12'sd-1037, 11'sd812, 13'sd2466}, {13'sd2780, 9'sd227, 11'sd-965}, {12'sd-1286, 11'sd628, 11'sd588}},
{{8'sd-104, 13'sd-2882, 13'sd-3004}, {12'sd-1380, 12'sd-1894, 13'sd-3298}, {11'sd790, 10'sd496, 12'sd-1765}},
{{12'sd2009, 12'sd-1542, 14'sd-4654}, {12'sd-1303, 12'sd1736, 5'sd15}, {14'sd4566, 10'sd-445, 12'sd1343}},
{{11'sd-979, 9'sd-203, 12'sd1800}, {12'sd-1308, 12'sd1128, 10'sd-333}, {13'sd-2383, 12'sd-1394, 10'sd256}},
{{13'sd-2383, 12'sd1999, 12'sd1835}, {13'sd2470, 10'sd-298, 12'sd-1718}, {13'sd2082, 11'sd990, 8'sd-112}},
{{13'sd-3119, 11'sd692, 12'sd-1248}, {7'sd50, 12'sd1565, 14'sd4483}, {11'sd677, 11'sd-556, 12'sd1170}},
{{13'sd2370, 11'sd-957, 11'sd-533}, {11'sd930, 11'sd-886, 13'sd-2931}, {11'sd951, 12'sd1271, 13'sd-3095}},
{{9'sd238, 10'sd-364, 13'sd-2471}, {9'sd-219, 13'sd-2899, 10'sd394}, {13'sd-2513, 11'sd-525, 13'sd2956}},
{{13'sd2975, 13'sd2429, 14'sd4485}, {13'sd-2184, 12'sd1215, 11'sd-884}, {12'sd-1474, 13'sd3636, 12'sd1503}},
{{11'sd-544, 13'sd-2440, 10'sd363}, {11'sd-673, 12'sd1695, 12'sd1105}, {10'sd-435, 11'sd575, 12'sd-1713}},
{{13'sd2158, 13'sd-2641, 11'sd868}, {13'sd-2326, 12'sd1234, 11'sd713}, {12'sd-1230, 4'sd-6, 13'sd2254}},
{{11'sd-560, 12'sd-1132, 13'sd2343}, {12'sd1332, 9'sd-201, 13'sd-2225}, {12'sd1103, 12'sd-2033, 10'sd-434}},
{{11'sd-890, 13'sd-2379, 12'sd-1515}, {9'sd218, 11'sd530, 12'sd1975}, {12'sd-1105, 12'sd-1602, 12'sd1675}},
{{11'sd-824, 11'sd-635, 13'sd2144}, {12'sd1818, 12'sd-1434, 12'sd1931}, {12'sd-1088, 10'sd427, 10'sd339}},
{{11'sd-586, 12'sd-1243, 13'sd-2276}, {12'sd-1478, 10'sd-433, 12'sd1661}, {13'sd2953, 11'sd-840, 11'sd-567}},
{{12'sd-1986, 13'sd-2768, 14'sd-5876}, {14'sd-4352, 12'sd1845, 14'sd-4563}, {11'sd753, 11'sd-981, 13'sd-4061}},
{{13'sd3178, 12'sd1967, 14'sd4559}, {12'sd2008, 11'sd-733, 13'sd2514}, {6'sd-20, 14'sd-4310, 11'sd-895}},
{{13'sd2732, 13'sd-2233, 13'sd-2774}, {13'sd-2626, 6'sd-30, 13'sd2347}, {11'sd-686, 13'sd-3159, 11'sd-758}},
{{13'sd2228, 13'sd-2515, 9'sd193}, {11'sd1016, 9'sd149, 13'sd2900}, {12'sd-1281, 11'sd-590, 12'sd-1305}},
{{10'sd382, 13'sd2240, 11'sd661}, {13'sd2376, 13'sd-2804, 12'sd-1959}, {13'sd-2095, 13'sd-2828, 12'sd-1613}},
{{12'sd-1353, 11'sd669, 10'sd256}, {13'sd2508, 11'sd-862, 10'sd498}, {13'sd-2964, 10'sd314, 13'sd2072}},
{{11'sd692, 12'sd-1188, 12'sd1405}, {12'sd1477, 10'sd-298, 12'sd1917}, {10'sd-389, 13'sd2136, 12'sd1262}},
{{13'sd2147, 13'sd3667, 12'sd1417}, {11'sd954, 12'sd1350, 13'sd-2980}, {12'sd1059, 10'sd263, 11'sd554}},
{{11'sd-532, 12'sd1706, 11'sd-805}, {12'sd1105, 12'sd-1712, 12'sd1202}, {13'sd2158, 10'sd337, 12'sd-1117}},
{{13'sd-3310, 9'sd-172, 14'sd-5385}, {12'sd-1451, 9'sd-218, 13'sd-2908}, {11'sd992, 13'sd2582, 10'sd-397}},
{{12'sd1805, 13'sd2325, 11'sd-908}, {11'sd-677, 13'sd-2063, 12'sd1146}, {14'sd-4635, 13'sd-3427, 13'sd2125}},
{{13'sd2751, 11'sd781, 12'sd1674}, {12'sd1219, 11'sd-944, 12'sd1125}, {12'sd-1991, 11'sd597, 12'sd-1988}},
{{10'sd-467, 10'sd305, 13'sd2847}, {12'sd-1631, 13'sd-2107, 12'sd-1520}, {12'sd-1622, 13'sd2729, 13'sd2940}},
{{13'sd2184, 11'sd-802, 12'sd1279}, {13'sd2934, 11'sd712, 13'sd-2457}, {13'sd3164, 13'sd-2351, 12'sd1245}},
{{14'sd4311, 11'sd715, 14'sd5094}, {12'sd-1449, 12'sd2000, 11'sd761}, {13'sd-4030, 12'sd-1785, 12'sd1620}},
{{11'sd778, 10'sd280, 12'sd1209}, {13'sd-2209, 10'sd-340, 13'sd-2068}, {11'sd693, 10'sd-407, 12'sd-1655}},
{{12'sd-1132, 11'sd699, 12'sd1554}, {13'sd-2742, 9'sd156, 13'sd2514}, {13'sd-2251, 12'sd1560, 9'sd-201}},
{{13'sd3291, 13'sd3022, 11'sd608}, {11'sd-1018, 10'sd502, 12'sd-1965}, {7'sd41, 11'sd1002, 14'sd-4502}},
{{10'sd-453, 13'sd2404, 12'sd1700}, {11'sd967, 12'sd-1486, 10'sd402}, {13'sd3610, 10'sd-465, 8'sd81}},
{{13'sd3728, 11'sd-736, 13'sd3827}, {13'sd3040, 11'sd-944, 13'sd4050}, {13'sd3122, 10'sd-294, 13'sd3170}},
{{11'sd1018, 12'sd1262, 11'sd613}, {12'sd-1864, 12'sd1734, 10'sd-406}, {12'sd-1724, 11'sd844, 12'sd1594}},
{{14'sd-4596, 12'sd-1528, 11'sd-1006}, {11'sd-954, 13'sd2635, 13'sd2344}, {10'sd411, 10'sd483, 12'sd1850}},
{{10'sd331, 13'sd3305, 12'sd1437}, {13'sd2070, 13'sd2171, 11'sd-557}, {13'sd-3807, 13'sd-2385, 13'sd2088}},
{{11'sd-834, 9'sd222, 12'sd-1074}, {13'sd2840, 12'sd1681, 6'sd-27}, {13'sd-2888, 13'sd2114, 11'sd-667}}},
{
{{10'sd455, 13'sd-2907, 12'sd-1734}, {11'sd1002, 12'sd1154, 13'sd-2178}, {12'sd1748, 7'sd39, 13'sd2783}},
{{13'sd-2562, 10'sd258, 12'sd1556}, {10'sd493, 12'sd-1782, 12'sd1996}, {12'sd-1642, 12'sd-1190, 13'sd-2411}},
{{11'sd-841, 12'sd1927, 11'sd818}, {13'sd2931, 13'sd-2216, 12'sd-1560}, {12'sd1493, 13'sd-2325, 12'sd1238}},
{{12'sd1373, 12'sd-1046, 12'sd1639}, {11'sd-869, 13'sd-2669, 9'sd-162}, {13'sd2118, 12'sd1516, 11'sd-594}},
{{12'sd1619, 12'sd1946, 10'sd355}, {10'sd-320, 12'sd1582, 12'sd1977}, {12'sd-1434, 12'sd-1959, 12'sd-1665}},
{{12'sd1392, 12'sd-1413, 11'sd-630}, {8'sd-114, 11'sd802, 12'sd1855}, {13'sd2461, 12'sd-1424, 11'sd822}},
{{10'sd-413, 13'sd2451, 13'sd2476}, {12'sd1096, 12'sd1386, 13'sd-2666}, {12'sd-1760, 12'sd2001, 11'sd535}},
{{12'sd-1180, 13'sd-2392, 13'sd-2553}, {12'sd1514, 10'sd494, 9'sd-224}, {13'sd2778, 13'sd2129, 12'sd-2027}},
{{9'sd-148, 12'sd-1118, 13'sd-2564}, {12'sd-2025, 13'sd-2599, 12'sd1238}, {13'sd3192, 13'sd2771, 5'sd-12}},
{{12'sd1723, 13'sd-2464, 12'sd-1530}, {13'sd2200, 12'sd-1096, 10'sd344}, {10'sd349, 10'sd297, 10'sd-343}},
{{12'sd1355, 13'sd2781, 12'sd-1997}, {13'sd2378, 12'sd-1070, 11'sd-867}, {12'sd1728, 5'sd-9, 12'sd1187}},
{{13'sd2351, 9'sd167, 8'sd-72}, {8'sd-106, 13'sd-2725, 12'sd-1100}, {12'sd-1464, 13'sd2514, 12'sd1940}},
{{12'sd1970, 12'sd-1834, 13'sd2514}, {13'sd-3032, 12'sd1142, 12'sd-1302}, {11'sd-906, 10'sd-492, 12'sd-1194}},
{{13'sd2722, 13'sd-2430, 10'sd493}, {9'sd-195, 13'sd-2601, 12'sd1148}, {13'sd-2407, 13'sd2051, 10'sd-461}},
{{13'sd-2336, 9'sd-252, 13'sd-2464}, {11'sd979, 12'sd1125, 13'sd-2147}, {12'sd-1277, 13'sd-2437, 10'sd285}},
{{11'sd623, 8'sd-101, 13'sd2636}, {11'sd519, 9'sd-173, 13'sd-2182}, {13'sd-2063, 12'sd1251, 12'sd1555}},
{{13'sd2877, 12'sd1313, 12'sd1834}, {12'sd1062, 9'sd218, 10'sd-380}, {8'sd79, 10'sd395, 13'sd-2257}},
{{12'sd-1420, 11'sd849, 10'sd273}, {12'sd1029, 9'sd-180, 13'sd2332}, {12'sd1321, 13'sd3050, 12'sd1284}},
{{11'sd-811, 12'sd-1435, 13'sd-3004}, {11'sd548, 9'sd-155, 11'sd-897}, {12'sd-1143, 13'sd-3098, 8'sd74}},
{{13'sd-2498, 11'sd-999, 13'sd2081}, {10'sd-377, 13'sd-2113, 12'sd1336}, {12'sd-2047, 12'sd-1089, 12'sd-1360}},
{{12'sd1156, 11'sd-668, 12'sd1697}, {12'sd-1223, 12'sd-1319, 13'sd-2586}, {13'sd3012, 11'sd539, 11'sd891}},
{{13'sd2363, 11'sd-809, 12'sd1598}, {13'sd-2643, 10'sd-389, 11'sd947}, {11'sd761, 12'sd-1149, 12'sd-1683}},
{{12'sd1105, 12'sd1114, 12'sd-1121}, {13'sd-2533, 12'sd1590, 12'sd1992}, {10'sd413, 8'sd-83, 13'sd-2440}},
{{12'sd1379, 12'sd-1103, 9'sd239}, {9'sd-183, 12'sd1705, 9'sd-139}, {12'sd-2025, 11'sd-562, 9'sd-174}},
{{12'sd-1289, 11'sd-672, 13'sd-2319}, {13'sd2213, 11'sd-563, 11'sd956}, {12'sd-1616, 7'sd-35, 7'sd-41}},
{{12'sd-1619, 10'sd393, 10'sd-267}, {10'sd266, 12'sd1469, 9'sd193}, {10'sd-361, 13'sd2400, 12'sd-1645}},
{{13'sd2332, 11'sd-832, 11'sd-525}, {12'sd-1083, 11'sd-669, 13'sd2215}, {13'sd-2189, 13'sd-3017, 12'sd-1292}},
{{13'sd2349, 8'sd80, 13'sd-2529}, {12'sd-1304, 12'sd-1974, 13'sd2283}, {12'sd1896, 13'sd-2257, 5'sd-15}},
{{9'sd151, 12'sd-1303, 7'sd-53}, {12'sd1915, 13'sd2283, 10'sd-326}, {13'sd-2576, 12'sd1093, 12'sd-1282}},
{{12'sd-1154, 10'sd399, 12'sd-1638}, {13'sd-2095, 13'sd-2431, 12'sd1519}, {12'sd-2045, 12'sd1831, 13'sd-2188}},
{{10'sd271, 13'sd2107, 11'sd-743}, {12'sd-1134, 11'sd612, 12'sd1993}, {11'sd-542, 13'sd-2811, 12'sd-1111}},
{{9'sd236, 11'sd-692, 6'sd26}, {11'sd-922, 10'sd439, 11'sd-585}, {13'sd2094, 9'sd-175, 12'sd1208}},
{{13'sd-2766, 9'sd231, 13'sd2577}, {10'sd-400, 9'sd161, 13'sd2240}, {12'sd1379, 13'sd-2339, 12'sd-1035}},
{{13'sd2058, 12'sd1921, 12'sd1196}, {13'sd-2220, 12'sd-1172, 12'sd-1714}, {10'sd380, 12'sd1173, 13'sd-2429}},
{{13'sd-2389, 12'sd1506, 12'sd-1273}, {13'sd2186, 12'sd1739, 11'sd868}, {13'sd2710, 12'sd2028, 11'sd662}},
{{11'sd-919, 10'sd472, 12'sd1538}, {11'sd-944, 12'sd-1933, 12'sd-1270}, {13'sd2326, 12'sd-1196, 12'sd-1120}},
{{11'sd982, 10'sd-497, 12'sd-1868}, {12'sd-1978, 11'sd1019, 11'sd-597}, {10'sd-462, 12'sd-1233, 13'sd-2237}},
{{13'sd-2164, 12'sd-1581, 13'sd2496}, {13'sd-2212, 11'sd-633, 10'sd465}, {11'sd-514, 12'sd1645, 10'sd408}},
{{11'sd688, 9'sd-252, 10'sd425}, {11'sd696, 11'sd-745, 12'sd-1055}, {11'sd941, 12'sd-1088, 10'sd409}},
{{13'sd-2579, 13'sd-2098, 11'sd519}, {12'sd1623, 11'sd-900, 13'sd-2659}, {12'sd-1520, 11'sd742, 12'sd1757}},
{{12'sd1370, 13'sd2432, 11'sd927}, {11'sd-628, 10'sd-427, 12'sd-1805}, {12'sd-1065, 12'sd-1277, 10'sd-290}},
{{11'sd-697, 12'sd1052, 12'sd1283}, {11'sd589, 10'sd432, 13'sd-2223}, {13'sd2304, 13'sd-2462, 11'sd757}},
{{10'sd458, 12'sd-1477, 12'sd1842}, {13'sd-2201, 12'sd-1149, 11'sd-565}, {12'sd1683, 12'sd-1699, 12'sd1363}},
{{13'sd2594, 10'sd-466, 12'sd-1446}, {13'sd-2056, 12'sd-1428, 10'sd-489}, {13'sd2523, 13'sd2674, 13'sd2922}},
{{10'sd423, 12'sd-1067, 13'sd-2077}, {12'sd1833, 11'sd625, 11'sd-612}, {9'sd-147, 11'sd-687, 10'sd350}},
{{10'sd272, 11'sd877, 12'sd-1337}, {12'sd1703, 12'sd-1214, 12'sd-1732}, {13'sd3065, 12'sd1108, 11'sd-577}},
{{12'sd1471, 13'sd-2372, 13'sd-2390}, {13'sd2825, 9'sd229, 12'sd1779}, {12'sd1226, 12'sd-1397, 11'sd-908}},
{{10'sd443, 12'sd-1134, 10'sd-507}, {11'sd891, 11'sd-711, 12'sd1404}, {11'sd-851, 11'sd-759, 13'sd-3089}},
{{9'sd-202, 12'sd-1449, 12'sd1533}, {13'sd-2509, 12'sd1053, 12'sd-1994}, {12'sd-1026, 12'sd-1105, 11'sd-715}},
{{12'sd1747, 8'sd64, 6'sd-23}, {11'sd825, 9'sd129, 11'sd611}, {12'sd-1943, 11'sd948, 13'sd2784}},
{{12'sd-1193, 13'sd2306, 13'sd-2264}, {13'sd2469, 12'sd-1599, 11'sd512}, {13'sd2707, 10'sd322, 13'sd-2830}},
{{11'sd-733, 12'sd1877, 12'sd-1395}, {11'sd785, 12'sd-1065, 12'sd-1998}, {13'sd-2648, 12'sd-1971, 11'sd-857}},
{{10'sd445, 13'sd-2271, 12'sd-1468}, {12'sd1559, 11'sd657, 9'sd-233}, {12'sd-1080, 11'sd967, 10'sd259}},
{{10'sd406, 13'sd-2391, 13'sd2415}, {12'sd-1149, 13'sd-2077, 12'sd-1849}, {13'sd-2817, 12'sd-1207, 12'sd-1725}},
{{11'sd871, 11'sd892, 12'sd1118}, {11'sd917, 13'sd-2733, 12'sd1241}, {12'sd-1547, 9'sd-129, 11'sd633}},
{{13'sd2156, 10'sd409, 13'sd-2360}, {11'sd567, 12'sd1912, 11'sd892}, {11'sd-956, 11'sd679, 11'sd-823}},
{{13'sd-2478, 13'sd-2590, 10'sd-323}, {12'sd-1491, 13'sd2581, 11'sd-560}, {13'sd-2710, 12'sd1348, 12'sd1474}},
{{11'sd964, 12'sd-1392, 12'sd-1395}, {12'sd1668, 12'sd-2000, 12'sd-1308}, {8'sd-83, 12'sd-2025, 11'sd557}},
{{12'sd1733, 9'sd-164, 13'sd2459}, {13'sd-2085, 12'sd-1762, 13'sd-2812}, {10'sd-388, 13'sd-2474, 9'sd-157}},
{{10'sd437, 13'sd2597, 13'sd-2263}, {12'sd2021, 12'sd1096, 12'sd-1479}, {12'sd-1130, 12'sd1453, 10'sd-292}},
{{12'sd-1582, 13'sd-2891, 13'sd-2163}, {12'sd1749, 12'sd1154, 13'sd-2822}, {13'sd-2381, 11'sd-656, 12'sd-1553}},
{{13'sd-2143, 12'sd1145, 9'sd-190}, {11'sd775, 12'sd-1747, 12'sd-1513}, {11'sd520, 12'sd-1756, 12'sd1555}},
{{9'sd246, 12'sd1557, 13'sd2237}, {12'sd1079, 13'sd-2318, 12'sd-1518}, {13'sd2146, 11'sd-726, 12'sd1279}},
{{13'sd2109, 10'sd-484, 12'sd2030}, {10'sd301, 11'sd-744, 9'sd-166}, {13'sd2441, 10'sd-356, 13'sd2350}}},
{
{{13'sd-2602, 12'sd1840, 13'sd2122}, {9'sd-231, 12'sd1208, 12'sd1883}, {12'sd-1267, 13'sd2372, 11'sd-873}},
{{13'sd-2356, 11'sd-744, 11'sd-681}, {12'sd-1843, 8'sd80, 13'sd-2639}, {12'sd2000, 12'sd-1530, 11'sd740}},
{{12'sd-1446, 12'sd-1846, 10'sd381}, {11'sd-540, 10'sd-386, 12'sd-1725}, {13'sd3100, 11'sd-661, 11'sd-641}},
{{10'sd-319, 10'sd-495, 11'sd749}, {13'sd2489, 12'sd1606, 12'sd-1620}, {8'sd114, 8'sd-111, 13'sd2254}},
{{11'sd670, 12'sd-1653, 12'sd-1341}, {13'sd-2227, 8'sd-71, 11'sd694}, {9'sd-137, 10'sd376, 11'sd-932}},
{{12'sd1623, 10'sd-456, 12'sd-1650}, {12'sd-1605, 13'sd-2254, 13'sd2489}, {11'sd858, 13'sd2386, 13'sd-2270}},
{{12'sd-1414, 12'sd1135, 12'sd-1330}, {12'sd1998, 13'sd2506, 11'sd560}, {13'sd2211, 9'sd-248, 11'sd-668}},
{{12'sd-1716, 12'sd-1785, 12'sd1316}, {10'sd-343, 13'sd2824, 12'sd-1785}, {9'sd-196, 13'sd-2326, 11'sd672}},
{{13'sd2225, 9'sd-252, 8'sd109}, {13'sd2646, 12'sd1293, 13'sd2419}, {12'sd-1711, 12'sd1716, 13'sd-2719}},
{{11'sd-862, 13'sd2768, 12'sd1707}, {6'sd26, 12'sd-1422, 12'sd-1147}, {12'sd-1347, 12'sd1059, 11'sd997}},
{{11'sd-859, 12'sd-1615, 13'sd-2687}, {13'sd-2482, 13'sd2087, 13'sd-2656}, {13'sd2118, 13'sd-2085, 10'sd265}},
{{12'sd1816, 13'sd-2078, 13'sd2633}, {13'sd-3006, 10'sd457, 12'sd1276}, {13'sd-2333, 12'sd-1397, 13'sd-2231}},
{{12'sd-1959, 13'sd4091, 13'sd2868}, {13'sd2583, 13'sd2934, 4'sd5}, {12'sd-1966, 11'sd849, 13'sd3952}},
{{12'sd1988, 10'sd-509, 11'sd882}, {10'sd-443, 12'sd-1856, 12'sd-1206}, {10'sd-420, 12'sd1508, 11'sd1009}},
{{13'sd-2519, 13'sd-2505, 11'sd-1023}, {11'sd-1019, 11'sd980, 11'sd-512}, {12'sd1459, 10'sd-431, 12'sd-1833}},
{{12'sd1185, 12'sd-1448, 11'sd-598}, {9'sd215, 10'sd342, 12'sd1413}, {12'sd1619, 12'sd1658, 10'sd-295}},
{{13'sd-2707, 12'sd-1816, 13'sd2371}, {13'sd2338, 11'sd-665, 11'sd-680}, {12'sd-1820, 11'sd-603, 12'sd1045}},
{{11'sd857, 6'sd-23, 12'sd-1481}, {6'sd-22, 12'sd-1540, 12'sd1241}, {13'sd2713, 12'sd-1811, 11'sd877}},
{{13'sd-2465, 13'sd-2480, 13'sd-2928}, {13'sd2206, 12'sd1408, 12'sd1668}, {13'sd-2076, 13'sd-2481, 13'sd-3476}},
{{13'sd-2427, 12'sd-1299, 11'sd668}, {12'sd1602, 12'sd1403, 13'sd-2104}, {11'sd783, 12'sd1814, 10'sd-373}},
{{13'sd2851, 7'sd-40, 13'sd-2810}, {13'sd2991, 12'sd-1028, 11'sd-684}, {13'sd2461, 12'sd-1333, 13'sd-2090}},
{{12'sd-1752, 12'sd1055, 13'sd2801}, {10'sd-312, 12'sd-1244, 9'sd-206}, {12'sd1482, 8'sd93, 9'sd-173}},
{{10'sd-474, 13'sd-2483, 12'sd-1380}, {13'sd2241, 9'sd-181, 11'sd980}, {12'sd1895, 10'sd323, 13'sd-2356}},
{{12'sd1926, 13'sd-3006, 10'sd-421}, {13'sd-2191, 10'sd-299, 12'sd-1256}, {13'sd2352, 12'sd1783, 8'sd-67}},
{{13'sd2748, 11'sd774, 12'sd-1340}, {13'sd2383, 10'sd505, 13'sd2395}, {12'sd1796, 12'sd-1450, 13'sd-2810}},
{{13'sd-2119, 13'sd-2564, 12'sd-1455}, {11'sd842, 11'sd-622, 12'sd1147}, {11'sd826, 13'sd-2805, 11'sd-879}},
{{11'sd890, 13'sd2418, 4'sd4}, {12'sd1949, 12'sd-1164, 13'sd3011}, {12'sd-1812, 12'sd1995, 12'sd-1290}},
{{12'sd-1632, 12'sd1424, 12'sd1248}, {11'sd734, 12'sd-1849, 13'sd2646}, {12'sd-1434, 11'sd-553, 11'sd647}},
{{12'sd-1742, 11'sd546, 9'sd229}, {12'sd1581, 12'sd1227, 12'sd2004}, {13'sd2720, 12'sd2024, 12'sd-1361}},
{{13'sd2432, 12'sd-1970, 11'sd-681}, {10'sd-443, 12'sd-1295, 13'sd2529}, {13'sd-2067, 11'sd974, 11'sd795}},
{{13'sd-2920, 13'sd-3108, 13'sd-3153}, {10'sd412, 12'sd-1397, 10'sd-395}, {12'sd1555, 13'sd-3659, 11'sd-895}},
{{11'sd-533, 11'sd-692, 13'sd2712}, {12'sd-1947, 12'sd-1256, 12'sd2006}, {10'sd442, 9'sd252, 12'sd1404}},
{{11'sd-1008, 13'sd-2987, 11'sd634}, {12'sd1946, 13'sd2211, 9'sd-255}, {13'sd-3058, 12'sd-1697, 9'sd243}},
{{12'sd-1471, 11'sd749, 10'sd301}, {12'sd1192, 12'sd1916, 9'sd177}, {13'sd-2508, 9'sd138, 12'sd-1793}},
{{11'sd962, 12'sd-1345, 12'sd-1650}, {13'sd-2360, 13'sd-2456, 11'sd-890}, {13'sd3026, 13'sd2146, 11'sd595}},
{{13'sd-2662, 11'sd-686, 12'sd-1747}, {12'sd-1270, 10'sd484, 12'sd1310}, {8'sd91, 11'sd624, 11'sd-806}},
{{12'sd1710, 12'sd1906, 12'sd-1840}, {11'sd696, 12'sd-1875, 13'sd2194}, {10'sd-385, 12'sd1790, 10'sd-464}},
{{11'sd-780, 11'sd975, 12'sd1769}, {13'sd-2343, 12'sd1934, 12'sd-1171}, {13'sd-2511, 13'sd2279, 12'sd1933}},
{{12'sd-2033, 13'sd-2486, 12'sd1921}, {12'sd-1998, 11'sd-918, 11'sd-663}, {8'sd65, 11'sd924, 12'sd-1235}},
{{12'sd-1425, 13'sd-2086, 13'sd2480}, {11'sd-828, 11'sd770, 10'sd438}, {9'sd-156, 13'sd2068, 12'sd-1631}},
{{11'sd685, 12'sd1906, 11'sd530}, {13'sd2461, 12'sd-1404, 12'sd1314}, {11'sd-593, 10'sd-408, 13'sd-2099}},
{{13'sd-2514, 13'sd2650, 13'sd2141}, {13'sd-2403, 11'sd897, 11'sd-827}, {13'sd2420, 12'sd-1604, 13'sd2883}},
{{13'sd2188, 13'sd2557, 10'sd491}, {13'sd2093, 12'sd-1077, 11'sd569}, {7'sd-63, 13'sd2386, 13'sd-2218}},
{{13'sd-2407, 11'sd578, 9'sd-232}, {12'sd-1505, 12'sd-1539, 11'sd848}, {11'sd-1016, 9'sd252, 13'sd2513}},
{{12'sd-1677, 13'sd2281, 12'sd-1621}, {11'sd-940, 13'sd3293, 11'sd898}, {12'sd1520, 13'sd3569, 12'sd-1406}},
{{13'sd-2617, 12'sd-1264, 10'sd373}, {13'sd-2183, 11'sd-590, 10'sd-430}, {13'sd-2121, 12'sd-1260, 12'sd1191}},
{{10'sd-393, 12'sd-1603, 8'sd-127}, {11'sd-905, 8'sd-93, 11'sd-935}, {12'sd2025, 12'sd-1555, 9'sd178}},
{{12'sd-1768, 10'sd375, 13'sd-2591}, {12'sd1103, 4'sd4, 12'sd1935}, {13'sd-3214, 12'sd1035, 9'sd142}},
{{12'sd1561, 13'sd-2285, 13'sd-2288}, {12'sd1967, 13'sd-2096, 12'sd1351}, {13'sd3034, 11'sd-955, 10'sd455}},
{{12'sd1076, 12'sd1699, 13'sd2750}, {11'sd724, 13'sd-2244, 11'sd-882}, {12'sd-1723, 10'sd444, 12'sd1633}},
{{13'sd-3584, 12'sd-1790, 8'sd-84}, {13'sd-2141, 13'sd2332, 12'sd-1356}, {13'sd-2342, 11'sd-577, 12'sd-1773}},
{{12'sd1720, 11'sd808, 12'sd-1668}, {12'sd1404, 12'sd1088, 12'sd-1710}, {12'sd1376, 9'sd-219, 13'sd2603}},
{{9'sd-251, 13'sd-2396, 10'sd461}, {11'sd1012, 8'sd-110, 11'sd-754}, {12'sd1667, 11'sd898, 12'sd-1495}},
{{8'sd87, 12'sd1713, 12'sd-1114}, {12'sd1203, 12'sd-1474, 13'sd-2531}, {13'sd2353, 12'sd-2013, 13'sd2353}},
{{13'sd-3267, 11'sd-941, 12'sd-1490}, {12'sd1552, 7'sd-58, 10'sd-275}, {12'sd-1882, 13'sd3222, 13'sd3094}},
{{11'sd585, 13'sd-2102, 12'sd1479}, {12'sd-1280, 13'sd-2275, 12'sd-1339}, {10'sd317, 10'sd434, 11'sd-699}},
{{13'sd-2853, 12'sd1293, 10'sd282}, {12'sd-1045, 13'sd-2177, 12'sd-1580}, {8'sd80, 13'sd2514, 13'sd2479}},
{{11'sd-588, 11'sd816, 13'sd-2116}, {12'sd1114, 12'sd1980, 12'sd2002}, {13'sd2944, 12'sd-1862, 12'sd1707}},
{{12'sd-1251, 13'sd2678, 12'sd1940}, {12'sd-1725, 12'sd1840, 13'sd2277}, {11'sd776, 11'sd592, 13'sd-2577}},
{{8'sd-126, 11'sd-873, 12'sd1305}, {13'sd-2882, 11'sd982, 11'sd952}, {12'sd-1616, 12'sd-1691, 10'sd-437}},
{{11'sd-1021, 9'sd-180, 12'sd-1129}, {11'sd1021, 13'sd-2339, 7'sd43}, {11'sd708, 11'sd528, 13'sd2110}},
{{11'sd707, 12'sd-1759, 13'sd2184}, {9'sd-136, 8'sd68, 11'sd636}, {11'sd-867, 11'sd-833, 12'sd-1617}},
{{12'sd-1332, 13'sd-2466, 11'sd932}, {11'sd-806, 11'sd-1018, 11'sd-1004}, {13'sd2741, 11'sd840, 10'sd-426}},
{{11'sd-910, 11'sd639, 11'sd613}, {11'sd-1007, 11'sd601, 13'sd-2876}, {11'sd847, 10'sd289, 12'sd-1801}}},
{
{{12'sd1878, 11'sd-951, 12'sd1106}, {13'sd2233, 11'sd-786, 13'sd2426}, {9'sd-132, 12'sd1718, 13'sd-2253}},
{{11'sd603, 9'sd-232, 11'sd900}, {11'sd-903, 9'sd-131, 12'sd1945}, {13'sd2795, 11'sd-596, 13'sd2553}},
{{12'sd1716, 11'sd-819, 12'sd1258}, {12'sd1117, 12'sd-1366, 13'sd2914}, {11'sd-693, 11'sd1015, 12'sd1446}},
{{11'sd-606, 12'sd-1650, 13'sd2469}, {12'sd-1431, 11'sd-516, 7'sd44}, {11'sd904, 12'sd-1465, 12'sd-1702}},
{{12'sd1597, 9'sd155, 13'sd-2145}, {11'sd758, 11'sd-808, 13'sd2309}, {11'sd723, 10'sd281, 13'sd-2233}},
{{12'sd-2024, 12'sd1214, 8'sd87}, {12'sd-1675, 12'sd1661, 13'sd-2395}, {9'sd-142, 12'sd1581, 11'sd876}},
{{12'sd1304, 13'sd-2709, 13'sd-2792}, {12'sd-1202, 13'sd-2353, 12'sd-1790}, {10'sd-441, 12'sd-1092, 6'sd29}},
{{13'sd2310, 11'sd773, 11'sd-702}, {9'sd142, 12'sd-1584, 13'sd2843}, {12'sd1319, 12'sd-1466, 13'sd-2394}},
{{13'sd-2543, 11'sd-862, 12'sd1066}, {13'sd-3072, 11'sd-936, 11'sd-892}, {11'sd704, 11'sd-696, 13'sd-2520}},
{{13'sd2247, 12'sd1567, 12'sd-1470}, {12'sd-1507, 13'sd2421, 12'sd-1957}, {13'sd2487, 11'sd1010, 11'sd850}},
{{12'sd-1761, 13'sd-2816, 12'sd-1485}, {12'sd1979, 12'sd-1055, 12'sd-1716}, {7'sd51, 12'sd-1259, 12'sd1767}},
{{9'sd199, 13'sd2456, 12'sd-1314}, {11'sd893, 10'sd-340, 13'sd2603}, {12'sd-1613, 11'sd-659, 9'sd-209}},
{{13'sd-2739, 12'sd-1843, 10'sd-297}, {12'sd-1897, 14'sd-4167, 12'sd-1230}, {10'sd-470, 8'sd117, 10'sd369}},
{{12'sd-1480, 12'sd1686, 13'sd2464}, {11'sd-750, 11'sd-959, 11'sd-736}, {13'sd2231, 12'sd-2006, 13'sd2471}},
{{12'sd-1457, 12'sd1443, 12'sd2028}, {10'sd454, 12'sd1090, 11'sd869}, {13'sd-2992, 13'sd2276, 12'sd1392}},
{{12'sd1293, 9'sd152, 8'sd76}, {10'sd-330, 13'sd2235, 12'sd-1709}, {13'sd-2671, 11'sd852, 12'sd-1456}},
{{13'sd-2100, 12'sd1652, 11'sd-1013}, {12'sd1711, 11'sd649, 13'sd2166}, {11'sd732, 10'sd-326, 13'sd3049}},
{{13'sd-3320, 12'sd1227, 10'sd298}, {12'sd1367, 11'sd799, 12'sd1991}, {11'sd898, 13'sd-2381, 13'sd-2608}},
{{10'sd-448, 12'sd-1088, 13'sd-2414}, {12'sd-1921, 12'sd-1496, 12'sd1258}, {13'sd2470, 9'sd-249, 12'sd1726}},
{{13'sd-2247, 12'sd1293, 13'sd-2072}, {12'sd1777, 13'sd-3101, 13'sd-2408}, {12'sd-1728, 11'sd715, 12'sd1571}},
{{11'sd689, 10'sd436, 13'sd2883}, {12'sd1122, 13'sd-2298, 13'sd2904}, {12'sd-2011, 12'sd-1888, 12'sd1369}},
{{11'sd-544, 11'sd863, 12'sd-1109}, {11'sd-862, 13'sd-2663, 12'sd-1748}, {13'sd-2282, 12'sd1754, 11'sd-742}},
{{10'sd309, 12'sd-1920, 13'sd-2218}, {9'sd-211, 11'sd515, 12'sd1962}, {8'sd-73, 12'sd-1883, 12'sd1296}},
{{13'sd-2050, 12'sd1788, 12'sd-1498}, {11'sd-593, 13'sd3193, 13'sd3188}, {8'sd-93, 12'sd1438, 9'sd182}},
{{12'sd-1545, 13'sd-2796, 10'sd-334}, {12'sd-1074, 13'sd-2108, 13'sd-2732}, {11'sd-921, 13'sd-2223, 13'sd2163}},
{{12'sd-1243, 13'sd-2149, 9'sd190}, {13'sd-2393, 12'sd-1342, 11'sd825}, {12'sd1156, 12'sd-1875, 13'sd-2142}},
{{11'sd556, 13'sd2971, 12'sd-1287}, {12'sd1343, 5'sd-11, 12'sd1976}, {9'sd-223, 12'sd1668, 12'sd1830}},
{{12'sd1118, 12'sd-1387, 11'sd-857}, {11'sd777, 12'sd-1694, 12'sd1534}, {13'sd3102, 13'sd3433, 12'sd-1420}},
{{13'sd2092, 11'sd-932, 12'sd-1582}, {13'sd-2836, 10'sd427, 10'sd260}, {11'sd-878, 10'sd365, 10'sd319}},
{{12'sd-1946, 13'sd2366, 12'sd-1923}, {11'sd739, 10'sd-506, 13'sd-2509}, {11'sd961, 12'sd-1797, 12'sd1758}},
{{10'sd436, 11'sd556, 13'sd-2184}, {10'sd-259, 12'sd-1475, 12'sd1652}, {13'sd3121, 7'sd-53, 12'sd1801}},
{{13'sd2726, 13'sd3113, 13'sd3257}, {10'sd351, 12'sd-1271, 12'sd-1578}, {12'sd1079, 12'sd2007, 10'sd-393}},
{{12'sd1355, 11'sd-670, 12'sd-1108}, {13'sd2350, 10'sd-335, 12'sd1218}, {13'sd2311, 13'sd2702, 12'sd1605}},
{{11'sd645, 13'sd2361, 12'sd1564}, {9'sd-251, 10'sd388, 12'sd-1267}, {12'sd1757, 12'sd1228, 8'sd-120}},
{{9'sd-225, 13'sd-2739, 11'sd681}, {13'sd-2280, 12'sd1140, 12'sd-1563}, {12'sd1883, 12'sd-1565, 11'sd-702}},
{{12'sd1367, 11'sd-1021, 11'sd802}, {13'sd-2207, 13'sd-2644, 13'sd-2529}, {8'sd-101, 12'sd1376, 12'sd-1650}},
{{12'sd-1615, 12'sd-1924, 12'sd1238}, {12'sd1122, 11'sd815, 12'sd1696}, {12'sd1577, 11'sd-892, 12'sd1523}},
{{12'sd-1437, 12'sd-1835, 11'sd-611}, {13'sd-2067, 13'sd-2068, 12'sd1132}, {13'sd2153, 13'sd-2149, 12'sd1493}},
{{13'sd2303, 12'sd1418, 12'sd-1422}, {12'sd-1768, 12'sd1368, 13'sd2540}, {12'sd1753, 13'sd-2812, 13'sd-2679}},
{{12'sd1720, 12'sd-1639, 8'sd-115}, {11'sd928, 12'sd-1101, 10'sd388}, {7'sd47, 13'sd2849, 12'sd1504}},
{{11'sd-1000, 10'sd-360, 11'sd864}, {12'sd-1873, 12'sd1090, 11'sd871}, {12'sd1357, 13'sd2400, 10'sd371}},
{{12'sd-1578, 11'sd-699, 12'sd-1823}, {11'sd809, 9'sd-206, 10'sd317}, {11'sd928, 10'sd507, 13'sd-3482}},
{{13'sd-2456, 12'sd-1861, 12'sd-1058}, {13'sd-2091, 12'sd1640, 10'sd-483}, {12'sd1389, 13'sd-2104, 11'sd-603}},
{{8'sd-111, 12'sd-1157, 10'sd-505}, {11'sd-1004, 12'sd1545, 7'sd57}, {13'sd-2454, 13'sd-2257, 13'sd-2071}},
{{12'sd-1483, 13'sd-2214, 11'sd802}, {13'sd2056, 11'sd846, 12'sd-2043}, {12'sd1985, 11'sd895, 11'sd930}},
{{10'sd403, 13'sd2064, 11'sd-903}, {13'sd-2521, 11'sd-894, 13'sd-2611}, {4'sd-5, 11'sd-874, 10'sd-304}},
{{13'sd-3029, 11'sd-922, 10'sd-451}, {8'sd-71, 11'sd720, 11'sd981}, {12'sd-1355, 13'sd-2171, 10'sd-329}},
{{13'sd3267, 11'sd-940, 11'sd767}, {11'sd760, 12'sd1759, 10'sd387}, {13'sd2298, 12'sd1876, 7'sd57}},
{{11'sd884, 12'sd-1851, 12'sd1142}, {13'sd-2409, 10'sd-296, 12'sd1966}, {12'sd-1700, 12'sd-1551, 13'sd3335}},
{{12'sd-1417, 10'sd455, 12'sd-1968}, {12'sd1514, 13'sd-2758, 10'sd-281}, {11'sd562, 12'sd-1180, 9'sd194}},
{{11'sd556, 12'sd-1396, 13'sd3481}, {13'sd3563, 13'sd2728, 11'sd588}, {10'sd341, 12'sd1203, 13'sd2194}},
{{13'sd-2081, 8'sd82, 12'sd1673}, {9'sd231, 13'sd-2179, 12'sd-1307}, {12'sd-1717, 11'sd-515, 12'sd-1783}},
{{13'sd-2586, 12'sd1171, 13'sd2492}, {11'sd-974, 11'sd856, 13'sd-2356}, {12'sd1327, 13'sd2390, 12'sd-1786}},
{{12'sd-1528, 11'sd949, 12'sd-1987}, {12'sd1621, 9'sd169, 11'sd665}, {12'sd-1682, 11'sd-974, 12'sd1782}},
{{13'sd2530, 12'sd1616, 12'sd1505}, {13'sd2620, 10'sd-468, 12'sd-1605}, {11'sd684, 11'sd-780, 13'sd-2608}},
{{13'sd-2871, 13'sd2112, 12'sd1524}, {12'sd1829, 12'sd1767, 11'sd-590}, {13'sd-2329, 12'sd1749, 13'sd-3231}},
{{12'sd1979, 13'sd3038, 11'sd589}, {9'sd128, 11'sd898, 11'sd549}, {11'sd762, 12'sd1844, 10'sd360}},
{{11'sd-849, 10'sd-426, 8'sd-82}, {9'sd221, 12'sd1114, 12'sd-1528}, {13'sd2976, 12'sd-1602, 13'sd2095}},
{{11'sd-822, 13'sd-2332, 12'sd-1987}, {12'sd-1511, 12'sd-1613, 13'sd-2136}, {13'sd2992, 13'sd2666, 12'sd-1139}},
{{12'sd-1103, 11'sd-789, 12'sd-1217}, {13'sd-2104, 12'sd2011, 10'sd-260}, {11'sd-730, 13'sd-3130, 12'sd-1416}},
{{13'sd2112, 12'sd1582, 11'sd779}, {13'sd2363, 10'sd295, 10'sd342}, {12'sd-2044, 12'sd1470, 12'sd-1674}},
{{11'sd979, 11'sd705, 9'sd-237}, {6'sd-31, 12'sd1355, 12'sd-1697}, {13'sd2398, 13'sd2241, 11'sd861}},
{{11'sd-803, 10'sd-262, 9'sd135}, {13'sd2392, 13'sd-2650, 11'sd-950}, {12'sd-1145, 12'sd1094, 12'sd1585}},
{{11'sd-883, 12'sd1090, 12'sd1729}, {12'sd-1619, 11'sd1010, 10'sd423}, {8'sd-74, 11'sd-564, 12'sd-1831}}},
{
{{11'sd-628, 12'sd-1887, 12'sd1132}, {11'sd-909, 11'sd-923, 11'sd-958}, {12'sd-1798, 13'sd2376, 12'sd-1858}},
{{12'sd-1962, 11'sd638, 12'sd1389}, {11'sd997, 11'sd-879, 12'sd-1175}, {13'sd2191, 12'sd1605, 10'sd-340}},
{{13'sd-2345, 13'sd-2585, 12'sd1626}, {13'sd2633, 13'sd2490, 12'sd-1228}, {13'sd-3124, 13'sd2056, 12'sd1191}},
{{12'sd-1041, 10'sd-404, 12'sd2016}, {12'sd-1737, 12'sd-1161, 13'sd2469}, {12'sd-1526, 12'sd-1275, 12'sd1257}},
{{12'sd-1821, 10'sd-324, 13'sd2553}, {13'sd-2097, 12'sd-1119, 11'sd672}, {13'sd2209, 12'sd1719, 13'sd2298}},
{{6'sd-26, 12'sd1852, 12'sd-1480}, {12'sd1770, 11'sd746, 13'sd-2327}, {13'sd2055, 12'sd1890, 12'sd-1402}},
{{10'sd335, 13'sd-2595, 7'sd60}, {13'sd2103, 11'sd704, 12'sd1986}, {13'sd3538, 11'sd999, 11'sd860}},
{{12'sd-1841, 12'sd1258, 13'sd-2109}, {13'sd2458, 12'sd1391, 13'sd2585}, {12'sd1458, 10'sd-325, 12'sd-1625}},
{{12'sd1191, 13'sd-2162, 10'sd397}, {12'sd-1684, 11'sd716, 12'sd1904}, {12'sd1935, 8'sd-122, 10'sd470}},
{{12'sd1775, 11'sd-708, 10'sd-437}, {13'sd-2221, 12'sd1733, 9'sd200}, {13'sd2764, 12'sd1854, 12'sd-1171}},
{{10'sd-309, 11'sd562, 13'sd-3144}, {13'sd-2387, 13'sd-2904, 12'sd-1916}, {10'sd-468, 11'sd-661, 13'sd2221}},
{{13'sd-2609, 13'sd2321, 13'sd-2522}, {9'sd212, 11'sd-876, 10'sd281}, {12'sd-1994, 13'sd2234, 12'sd-1136}},
{{13'sd-2455, 12'sd1589, 11'sd-711}, {12'sd1680, 10'sd264, 13'sd2395}, {12'sd1058, 13'sd3131, 13'sd3387}},
{{13'sd-2191, 13'sd-2725, 11'sd-636}, {13'sd2545, 9'sd250, 11'sd-792}, {9'sd220, 11'sd659, 8'sd-64}},
{{6'sd-29, 13'sd-2530, 12'sd1529}, {11'sd545, 13'sd2817, 11'sd801}, {12'sd-1220, 13'sd2085, 10'sd464}},
{{13'sd2525, 12'sd1697, 7'sd-34}, {10'sd335, 11'sd-658, 10'sd-479}, {11'sd-780, 11'sd-802, 7'sd-49}},
{{9'sd162, 12'sd-1454, 11'sd575}, {10'sd457, 12'sd1412, 10'sd-492}, {13'sd2640, 13'sd2079, 12'sd1133}},
{{11'sd686, 10'sd259, 13'sd-2862}, {12'sd1466, 12'sd1828, 11'sd-872}, {12'sd1905, 12'sd1913, 13'sd2288}},
{{11'sd-826, 12'sd1769, 12'sd1982}, {12'sd-1805, 13'sd-2084, 13'sd2939}, {11'sd-719, 12'sd1278, 11'sd652}},
{{13'sd-2820, 10'sd-414, 6'sd-16}, {12'sd-1489, 12'sd-1530, 13'sd2058}, {10'sd336, 12'sd1128, 13'sd-2740}},
{{11'sd572, 13'sd2441, 12'sd-1568}, {10'sd425, 11'sd951, 13'sd-2343}, {12'sd-1651, 12'sd1873, 11'sd868}},
{{12'sd-1837, 13'sd2199, 12'sd1995}, {12'sd-1130, 12'sd1236, 12'sd1041}, {13'sd3264, 13'sd2746, 13'sd2049}},
{{9'sd-206, 12'sd1687, 12'sd-1883}, {13'sd2060, 13'sd2049, 13'sd2165}, {13'sd2314, 12'sd-1541, 12'sd-1133}},
{{12'sd1616, 11'sd-848, 13'sd2743}, {12'sd1898, 11'sd-717, 11'sd-1013}, {13'sd2586, 12'sd1900, 10'sd325}},
{{11'sd-938, 11'sd-983, 10'sd300}, {10'sd-365, 12'sd1673, 7'sd-40}, {12'sd-1925, 13'sd-2791, 13'sd-2889}},
{{12'sd-1223, 12'sd1570, 13'sd-2617}, {11'sd568, 12'sd1706, 11'sd856}, {13'sd2473, 12'sd1200, 13'sd-2484}},
{{9'sd245, 9'sd153, 12'sd1987}, {13'sd2718, 10'sd329, 12'sd1250}, {9'sd-142, 12'sd-1109, 13'sd3111}},
{{12'sd-1686, 12'sd-1614, 12'sd1036}, {12'sd-1914, 12'sd-1466, 12'sd-1464}, {12'sd-1954, 13'sd2688, 12'sd-1087}},
{{11'sd-768, 12'sd-1115, 13'sd-2345}, {13'sd2260, 12'sd-1957, 13'sd2508}, {12'sd2012, 11'sd-548, 12'sd1989}},
{{12'sd1595, 10'sd501, 12'sd1267}, {13'sd-2849, 12'sd1271, 7'sd-49}, {13'sd-2073, 12'sd2028, 7'sd-56}},
{{12'sd-1499, 13'sd-2717, 9'sd171}, {13'sd2086, 11'sd-860, 13'sd-4039}, {13'sd2726, 12'sd-1656, 10'sd316}},
{{13'sd2773, 9'sd170, 10'sd332}, {11'sd954, 11'sd648, 12'sd1922}, {11'sd903, 13'sd2746, 12'sd-1761}},
{{9'sd-176, 11'sd582, 12'sd1220}, {13'sd2809, 12'sd-1630, 9'sd232}, {9'sd-245, 10'sd-392, 11'sd732}},
{{13'sd-2077, 9'sd-183, 12'sd-1591}, {12'sd1811, 13'sd-2427, 12'sd-1566}, {13'sd-2239, 13'sd-2711, 13'sd-3169}},
{{10'sd362, 12'sd1974, 12'sd1522}, {11'sd939, 11'sd-682, 11'sd917}, {8'sd87, 12'sd1682, 12'sd1280}},
{{12'sd-1793, 10'sd393, 11'sd646}, {10'sd500, 12'sd-1555, 11'sd-601}, {9'sd-165, 13'sd-2832, 12'sd-1926}},
{{13'sd2532, 11'sd-890, 13'sd2852}, {12'sd1983, 12'sd-1946, 13'sd2558}, {12'sd-1989, 12'sd1875, 12'sd1167}},
{{13'sd-2913, 11'sd683, 13'sd-2242}, {12'sd-1872, 4'sd-7, 11'sd674}, {12'sd1734, 10'sd382, 12'sd1521}},
{{13'sd2300, 12'sd1729, 11'sd-747}, {13'sd-2572, 12'sd1324, 8'sd-116}, {11'sd835, 12'sd-2006, 12'sd-1831}},
{{8'sd-71, 12'sd-1198, 9'sd198}, {11'sd-825, 11'sd551, 13'sd-2314}, {12'sd-1270, 13'sd2072, 11'sd-701}},
{{11'sd-711, 10'sd290, 12'sd1149}, {12'sd1732, 10'sd346, 12'sd-1474}, {13'sd3008, 11'sd-699, 12'sd1118}},
{{11'sd791, 13'sd-2139, 11'sd776}, {13'sd-2571, 10'sd291, 12'sd-1441}, {13'sd2276, 13'sd-2083, 12'sd-1993}},
{{11'sd574, 12'sd1405, 10'sd295}, {10'sd476, 13'sd-2299, 13'sd-2128}, {13'sd2481, 10'sd-404, 9'sd-156}},
{{13'sd-2971, 12'sd1884, 11'sd-791}, {9'sd195, 9'sd-188, 12'sd-1070}, {8'sd-96, 12'sd1918, 13'sd2409}},
{{12'sd-1689, 13'sd2297, 11'sd715}, {13'sd-2544, 12'sd1640, 11'sd-855}, {12'sd1145, 12'sd-1783, 10'sd-275}},
{{13'sd-2369, 12'sd-1864, 12'sd1867}, {9'sd-155, 10'sd-440, 10'sd-294}, {13'sd-2142, 10'sd369, 12'sd1418}},
{{11'sd-827, 13'sd2186, 12'sd1280}, {12'sd-1962, 10'sd-315, 13'sd-2945}, {11'sd-881, 12'sd-1538, 12'sd-1897}},
{{11'sd900, 12'sd-1723, 11'sd-776}, {12'sd-1622, 13'sd2308, 13'sd-2190}, {9'sd169, 13'sd3580, 13'sd-2178}},
{{10'sd434, 10'sd-428, 13'sd-2665}, {12'sd-1508, 12'sd2035, 12'sd-1486}, {11'sd-828, 13'sd-2336, 12'sd-1138}},
{{6'sd-26, 13'sd3088, 12'sd-1233}, {13'sd2553, 10'sd-281, 13'sd2082}, {11'sd-909, 7'sd42, 13'sd2878}},
{{12'sd-1530, 11'sd-863, 10'sd451}, {12'sd1663, 13'sd-2081, 12'sd1412}, {13'sd-2313, 12'sd-1236, 13'sd2913}},
{{13'sd2604, 12'sd1708, 13'sd-2769}, {10'sd371, 10'sd-331, 12'sd-1722}, {12'sd1626, 10'sd301, 12'sd-1530}},
{{12'sd1427, 12'sd1172, 13'sd2275}, {13'sd2147, 13'sd-2439, 7'sd37}, {12'sd1789, 10'sd298, 12'sd1629}},
{{13'sd2565, 11'sd-627, 12'sd1612}, {12'sd-1954, 13'sd-2316, 13'sd2358}, {13'sd-2492, 12'sd1134, 13'sd2549}},
{{12'sd-1266, 8'sd-118, 9'sd-238}, {8'sd-123, 12'sd-1976, 13'sd-2574}, {13'sd3425, 11'sd705, 11'sd617}},
{{4'sd-6, 11'sd857, 12'sd-1160}, {12'sd-1651, 13'sd-2118, 13'sd2495}, {11'sd923, 6'sd-25, 12'sd1061}},
{{13'sd2795, 6'sd25, 12'sd1684}, {13'sd-2178, 11'sd-780, 6'sd-26}, {11'sd923, 12'sd1336, 12'sd-1682}},
{{12'sd-1200, 12'sd1225, 10'sd286}, {9'sd225, 12'sd2011, 12'sd-1396}, {11'sd970, 13'sd2214, 11'sd-650}},
{{9'sd-145, 13'sd-2402, 13'sd2175}, {10'sd-261, 8'sd88, 9'sd-158}, {7'sd56, 11'sd960, 10'sd-475}},
{{13'sd-2703, 9'sd217, 12'sd-1804}, {12'sd1690, 12'sd1610, 13'sd2699}, {12'sd1256, 7'sd-59, 13'sd-2745}},
{{12'sd-1877, 12'sd1858, 12'sd-1724}, {12'sd-1230, 11'sd981, 11'sd-615}, {13'sd-2442, 12'sd-1604, 12'sd1210}},
{{12'sd-1350, 12'sd-1880, 13'sd2226}, {12'sd-1280, 9'sd-173, 12'sd1636}, {13'sd3130, 12'sd1082, 12'sd1650}},
{{11'sd858, 9'sd160, 12'sd-1046}, {11'sd778, 13'sd-2223, 12'sd1963}, {13'sd-2458, 12'sd-1572, 10'sd-481}},
{{12'sd1971, 12'sd1691, 11'sd978}, {13'sd-2695, 13'sd-2615, 13'sd-2539}, {12'sd1178, 13'sd2148, 12'sd1037}}},
{
{{13'sd2151, 11'sd810, 12'sd1383}, {12'sd1740, 13'sd-2877, 12'sd1313}, {13'sd-3174, 12'sd1424, 10'sd417}},
{{12'sd-1594, 12'sd-1911, 10'sd487}, {12'sd-1833, 8'sd-103, 9'sd219}, {10'sd508, 12'sd-1597, 13'sd2214}},
{{13'sd2396, 12'sd-1784, 10'sd-294}, {12'sd-1640, 11'sd629, 7'sd-43}, {11'sd-761, 12'sd1851, 12'sd-1201}},
{{10'sd-385, 9'sd-142, 8'sd104}, {13'sd3005, 11'sd-993, 12'sd1718}, {12'sd-1364, 8'sd74, 12'sd1634}},
{{12'sd1491, 13'sd2282, 12'sd-1589}, {11'sd988, 13'sd2497, 13'sd-2056}, {12'sd1971, 12'sd-1460, 9'sd-162}},
{{11'sd-951, 11'sd-573, 13'sd-2235}, {12'sd-1791, 12'sd1736, 12'sd1618}, {12'sd-1293, 12'sd1352, 11'sd-880}},
{{12'sd-1659, 13'sd-2224, 11'sd-801}, {11'sd961, 13'sd2320, 12'sd1992}, {11'sd950, 11'sd-770, 11'sd-947}},
{{12'sd1679, 11'sd-995, 13'sd-2842}, {13'sd2532, 12'sd1176, 12'sd-1537}, {12'sd-1894, 13'sd2936, 11'sd580}},
{{11'sd-643, 13'sd3275, 12'sd1127}, {13'sd2776, 13'sd3441, 12'sd-1706}, {9'sd202, 10'sd369, 12'sd1394}},
{{13'sd-2327, 11'sd-786, 11'sd528}, {11'sd-533, 12'sd1051, 12'sd-1228}, {12'sd1744, 10'sd481, 10'sd398}},
{{10'sd304, 12'sd1137, 8'sd-107}, {12'sd-1218, 13'sd2158, 13'sd2120}, {12'sd1205, 13'sd2450, 12'sd1795}},
{{12'sd-1087, 10'sd448, 10'sd-260}, {11'sd959, 12'sd-1347, 13'sd2289}, {10'sd-454, 12'sd1924, 12'sd-1070}},
{{13'sd-2260, 12'sd1326, 12'sd1491}, {12'sd-1031, 10'sd353, 13'sd2189}, {13'sd3304, 12'sd1884, 13'sd3339}},
{{12'sd1291, 10'sd-286, 11'sd-884}, {12'sd-1640, 11'sd-515, 12'sd1886}, {12'sd1533, 13'sd2527, 12'sd-1356}},
{{12'sd1806, 10'sd297, 13'sd2542}, {11'sd781, 8'sd-110, 11'sd632}, {12'sd-1697, 10'sd346, 11'sd-564}},
{{13'sd-2214, 13'sd-2766, 13'sd2071}, {13'sd-2496, 12'sd1477, 9'sd-228}, {7'sd48, 13'sd2174, 12'sd1892}},
{{13'sd2561, 13'sd-2293, 11'sd863}, {12'sd-1722, 13'sd2056, 11'sd991}, {11'sd-907, 12'sd-1401, 11'sd666}},
{{10'sd373, 10'sd377, 13'sd-3701}, {10'sd-424, 12'sd1612, 13'sd-2841}, {13'sd2962, 11'sd-516, 12'sd1662}},
{{13'sd-2325, 13'sd-2172, 10'sd372}, {12'sd-1460, 12'sd1544, 8'sd-93}, {12'sd-1887, 13'sd2242, 12'sd-1358}},
{{10'sd384, 12'sd-1258, 12'sd-1861}, {12'sd1578, 12'sd-1521, 11'sd827}, {11'sd-836, 11'sd-591, 13'sd-2251}},
{{11'sd-693, 13'sd2600, 12'sd1231}, {12'sd2041, 8'sd-102, 12'sd1269}, {13'sd-2415, 11'sd-746, 12'sd-1323}},
{{13'sd-2259, 13'sd-2239, 10'sd496}, {13'sd-2137, 12'sd-1127, 13'sd2101}, {12'sd1276, 10'sd349, 12'sd1484}},
{{13'sd-2510, 12'sd-1217, 13'sd-2127}, {13'sd3085, 13'sd-2232, 12'sd-1283}, {11'sd866, 13'sd2483, 11'sd541}},
{{12'sd1434, 11'sd-655, 12'sd1282}, {11'sd783, 12'sd-1346, 12'sd-1582}, {7'sd35, 10'sd480, 10'sd-472}},
{{11'sd-614, 12'sd-1427, 10'sd-334}, {11'sd-579, 10'sd484, 11'sd826}, {11'sd-955, 13'sd2315, 13'sd-2386}},
{{13'sd-2755, 12'sd1510, 12'sd2023}, {10'sd457, 13'sd2138, 12'sd1977}, {12'sd1215, 12'sd-1090, 12'sd-1796}},
{{12'sd1970, 11'sd-823, 11'sd543}, {11'sd-947, 13'sd3277, 13'sd2283}, {10'sd481, 12'sd-2030, 8'sd-98}},
{{12'sd1660, 12'sd-1909, 8'sd109}, {13'sd-2205, 13'sd-2089, 10'sd-413}, {12'sd-1076, 12'sd-1980, 12'sd-1319}},
{{13'sd-2063, 11'sd796, 10'sd493}, {13'sd-2347, 12'sd-1555, 13'sd-2498}, {13'sd-2544, 12'sd-1069, 12'sd-1219}},
{{12'sd1345, 11'sd-758, 11'sd-744}, {13'sd-2547, 13'sd-2529, 12'sd-1784}, {13'sd-2571, 13'sd-2897, 8'sd79}},
{{13'sd-3312, 10'sd-314, 13'sd-2457}, {11'sd-548, 10'sd370, 10'sd275}, {13'sd3696, 10'sd-437, 12'sd-1665}},
{{10'sd-386, 11'sd930, 13'sd2552}, {11'sd828, 13'sd-2296, 8'sd110}, {12'sd1627, 13'sd2062, 11'sd-903}},
{{10'sd312, 12'sd-1731, 11'sd-722}, {12'sd1782, 12'sd1254, 11'sd-546}, {10'sd370, 11'sd773, 13'sd-3544}},
{{12'sd-2044, 10'sd-289, 11'sd847}, {10'sd314, 12'sd-1768, 12'sd-1611}, {13'sd3138, 13'sd-3067, 8'sd96}},
{{10'sd494, 11'sd-606, 10'sd-373}, {13'sd-2489, 12'sd-1802, 13'sd-2581}, {11'sd993, 13'sd-2261, 12'sd-1993}},
{{10'sd275, 12'sd1191, 12'sd-1281}, {10'sd419, 10'sd418, 12'sd1184}, {11'sd-847, 12'sd-1426, 12'sd-1789}},
{{7'sd60, 13'sd2336, 12'sd1804}, {11'sd999, 13'sd-2460, 9'sd213}, {11'sd-888, 10'sd-286, 11'sd528}},
{{12'sd-1184, 13'sd-2420, 11'sd905}, {10'sd-438, 13'sd-2576, 11'sd828}, {12'sd-1378, 10'sd506, 8'sd112}},
{{10'sd-488, 9'sd140, 12'sd-1537}, {10'sd-311, 10'sd-350, 12'sd1714}, {10'sd-393, 12'sd-1714, 8'sd110}},
{{13'sd2241, 12'sd1940, 12'sd-1533}, {12'sd-1444, 11'sd612, 13'sd2066}, {9'sd209, 12'sd-1120, 11'sd870}},
{{11'sd-884, 10'sd-422, 12'sd-1965}, {12'sd-1349, 12'sd1191, 12'sd-1980}, {12'sd1371, 13'sd2292, 12'sd2005}},
{{12'sd1849, 9'sd142, 13'sd-2630}, {13'sd2402, 11'sd951, 13'sd2249}, {13'sd2486, 12'sd-1742, 13'sd2873}},
{{11'sd-629, 12'sd1693, 10'sd-322}, {12'sd1724, 13'sd2959, 13'sd-2089}, {12'sd1670, 12'sd1469, 13'sd2257}},
{{12'sd1647, 13'sd2270, 13'sd-2297}, {11'sd-741, 11'sd553, 9'sd-150}, {13'sd2326, 13'sd-2148, 13'sd2524}},
{{13'sd-2986, 13'sd2509, 9'sd171}, {12'sd1828, 13'sd2178, 12'sd1760}, {12'sd-1472, 12'sd1129, 9'sd-165}},
{{13'sd2253, 12'sd1486, 12'sd1519}, {10'sd-287, 13'sd2077, 13'sd-2288}, {12'sd1822, 12'sd1782, 12'sd-1384}},
{{11'sd580, 12'sd1271, 11'sd837}, {13'sd-2321, 12'sd-1793, 13'sd-2221}, {12'sd1636, 12'sd1674, 13'sd2165}},
{{13'sd-3757, 10'sd-476, 13'sd-2910}, {13'sd-3069, 13'sd-2311, 13'sd2510}, {11'sd757, 13'sd2164, 12'sd-1096}},
{{11'sd-761, 13'sd-3219, 10'sd388}, {10'sd293, 13'sd-2226, 13'sd-2361}, {10'sd440, 12'sd1400, 11'sd-607}},
{{8'sd80, 12'sd1524, 10'sd281}, {11'sd787, 10'sd256, 12'sd1213}, {12'sd-1675, 12'sd-1233, 13'sd-3644}},
{{13'sd-3861, 12'sd1421, 13'sd-2569}, {10'sd-261, 13'sd-2907, 11'sd809}, {10'sd281, 12'sd-1289, 13'sd-2252}},
{{11'sd-828, 12'sd1525, 12'sd-1900}, {11'sd-742, 13'sd2478, 11'sd-536}, {13'sd-2154, 11'sd875, 11'sd-787}},
{{12'sd1472, 12'sd-2029, 13'sd-2508}, {13'sd-2188, 12'sd1495, 12'sd-1543}, {13'sd2358, 12'sd1619, 12'sd1341}},
{{10'sd275, 11'sd841, 11'sd725}, {11'sd953, 13'sd3218, 12'sd1730}, {11'sd-779, 5'sd13, 12'sd-1429}},
{{13'sd-2239, 13'sd-2244, 12'sd-1487}, {13'sd-2362, 10'sd-509, 11'sd-688}, {12'sd1998, 11'sd-692, 12'sd1571}},
{{12'sd1539, 12'sd1032, 11'sd670}, {11'sd-836, 11'sd672, 12'sd-2000}, {13'sd-2529, 12'sd-1094, 12'sd1181}},
{{12'sd1454, 10'sd-418, 11'sd-882}, {13'sd-3350, 12'sd1849, 12'sd-1772}, {9'sd-130, 12'sd1094, 12'sd1964}},
{{11'sd619, 11'sd800, 12'sd1949}, {11'sd601, 12'sd1938, 13'sd2408}, {13'sd2321, 12'sd1599, 4'sd-5}},
{{13'sd2313, 10'sd-499, 11'sd-672}, {10'sd427, 13'sd-2253, 13'sd-2344}, {10'sd300, 11'sd737, 13'sd-2181}},
{{12'sd-1290, 10'sd256, 11'sd1012}, {13'sd2221, 12'sd-1671, 12'sd1689}, {12'sd2026, 11'sd799, 12'sd-1194}},
{{11'sd891, 12'sd1398, 12'sd-1286}, {10'sd-414, 13'sd-2554, 11'sd791}, {13'sd-2265, 13'sd2485, 12'sd-1100}},
{{12'sd-1336, 11'sd645, 12'sd-1910}, {12'sd-1726, 11'sd634, 12'sd-1566}, {13'sd2496, 9'sd-236, 11'sd771}},
{{13'sd-3136, 10'sd310, 12'sd1396}, {11'sd-704, 13'sd-2308, 13'sd-2242}, {13'sd2544, 11'sd825, 12'sd1454}},
{{12'sd-1656, 9'sd142, 13'sd-3083}, {13'sd-2182, 13'sd-2177, 12'sd1690}, {12'sd-1274, 11'sd1004, 11'sd-697}}},
{
{{12'sd1371, 12'sd-1287, 12'sd-1043}, {9'sd-245, 10'sd-399, 9'sd160}, {13'sd-3373, 13'sd-2670, 12'sd-1419}},
{{12'sd1919, 13'sd-2140, 12'sd1744}, {13'sd2268, 13'sd2247, 13'sd2150}, {13'sd2198, 12'sd-1816, 12'sd1374}},
{{10'sd360, 13'sd3996, 12'sd1128}, {12'sd1158, 10'sd-424, 12'sd1144}, {13'sd-2734, 12'sd1390, 12'sd-1636}},
{{10'sd-393, 12'sd-1750, 13'sd2847}, {12'sd1666, 11'sd813, 12'sd-1716}, {11'sd662, 13'sd-2878, 11'sd574}},
{{12'sd1390, 12'sd1970, 9'sd139}, {12'sd1424, 6'sd-26, 9'sd224}, {10'sd381, 11'sd-640, 12'sd-2016}},
{{11'sd-975, 13'sd-2434, 12'sd1551}, {13'sd-2365, 10'sd-330, 12'sd1087}, {13'sd2736, 11'sd889, 10'sd299}},
{{13'sd2416, 12'sd-1521, 13'sd3522}, {12'sd-1274, 13'sd-2783, 10'sd413}, {13'sd2148, 12'sd1677, 12'sd1383}},
{{11'sd-660, 11'sd822, 13'sd-2841}, {13'sd-2767, 13'sd2264, 12'sd-1249}, {12'sd-1239, 12'sd1039, 10'sd-282}},
{{13'sd-2899, 9'sd-213, 12'sd1429}, {11'sd-949, 12'sd-1195, 8'sd-121}, {13'sd2610, 10'sd277, 13'sd-2688}},
{{10'sd432, 12'sd1381, 12'sd1090}, {11'sd-577, 11'sd-569, 8'sd92}, {13'sd-2576, 13'sd2504, 11'sd825}},
{{10'sd-439, 12'sd2011, 12'sd1103}, {13'sd-2150, 9'sd-145, 11'sd1014}, {10'sd268, 10'sd279, 12'sd1831}},
{{12'sd1083, 9'sd-217, 12'sd1598}, {12'sd2025, 11'sd-866, 11'sd674}, {12'sd-1953, 11'sd-586, 8'sd76}},
{{13'sd2671, 7'sd-32, 12'sd-1182}, {13'sd-3271, 14'sd-4607, 11'sd-1001}, {11'sd657, 14'sd-5389, 14'sd-4359}},
{{10'sd-279, 12'sd-1890, 10'sd-262}, {10'sd351, 12'sd2039, 11'sd-861}, {10'sd390, 7'sd60, 13'sd-2785}},
{{11'sd-1005, 12'sd1212, 13'sd-2136}, {10'sd-340, 13'sd-2377, 12'sd-1029}, {12'sd1472, 11'sd620, 13'sd2588}},
{{11'sd-956, 10'sd395, 13'sd2048}, {12'sd1293, 6'sd-23, 13'sd2330}, {11'sd977, 12'sd1330, 13'sd-2244}},
{{13'sd2301, 13'sd2383, 13'sd2363}, {12'sd-1357, 12'sd-1272, 13'sd-2116}, {11'sd904, 13'sd-2144, 11'sd-980}},
{{9'sd143, 12'sd1915, 13'sd-3906}, {11'sd645, 12'sd-1342, 10'sd491}, {7'sd61, 12'sd1525, 11'sd-847}},
{{12'sd-1370, 12'sd-1036, 11'sd-824}, {11'sd583, 12'sd-1610, 10'sd-463}, {11'sd-679, 13'sd3298, 11'sd-815}},
{{11'sd-785, 13'sd2157, 10'sd-475}, {11'sd-925, 11'sd-747, 11'sd531}, {13'sd2268, 12'sd1313, 13'sd2353}},
{{12'sd1888, 11'sd617, 4'sd4}, {12'sd-1701, 11'sd1017, 11'sd695}, {12'sd-1814, 12'sd1064, 12'sd-1116}},
{{12'sd1620, 13'sd-2548, 13'sd2319}, {10'sd-445, 12'sd1164, 13'sd-2201}, {13'sd2167, 11'sd769, 12'sd1250}},
{{11'sd755, 13'sd2567, 13'sd-2070}, {12'sd1538, 11'sd530, 12'sd-1151}, {12'sd1570, 13'sd2383, 8'sd-95}},
{{8'sd110, 12'sd-1483, 13'sd-2709}, {12'sd1990, 13'sd-2143, 12'sd-1117}, {13'sd2548, 13'sd2418, 13'sd2489}},
{{13'sd2393, 13'sd-2315, 11'sd-619}, {12'sd-1690, 13'sd-2726, 11'sd724}, {8'sd-74, 11'sd909, 9'sd253}},
{{12'sd-1712, 11'sd-708, 10'sd471}, {12'sd-1860, 11'sd-820, 9'sd250}, {12'sd1358, 12'sd-1629, 12'sd1166}},
{{12'sd-1144, 10'sd-384, 12'sd1953}, {12'sd1372, 10'sd511, 9'sd-216}, {11'sd904, 11'sd-794, 9'sd224}},
{{13'sd2756, 12'sd-1067, 10'sd505}, {12'sd-1824, 10'sd463, 12'sd-1898}, {12'sd1905, 7'sd-45, 12'sd-1988}},
{{12'sd-1961, 8'sd-98, 13'sd3398}, {11'sd-785, 12'sd1587, 11'sd-968}, {12'sd-1451, 9'sd-255, 9'sd175}},
{{13'sd-2307, 12'sd1076, 12'sd-1445}, {12'sd-1559, 10'sd-461, 10'sd290}, {12'sd-1339, 9'sd224, 12'sd1339}},
{{13'sd-3649, 13'sd2437, 10'sd503}, {12'sd1819, 12'sd1654, 13'sd3089}, {13'sd2341, 12'sd1750, 12'sd1700}},
{{13'sd-2424, 12'sd1984, 11'sd-842}, {8'sd65, 13'sd-2167, 12'sd-1337}, {12'sd-1458, 12'sd-1054, 12'sd1688}},
{{12'sd-1325, 13'sd-2209, 13'sd-2558}, {12'sd-1357, 13'sd2513, 13'sd2104}, {10'sd-308, 13'sd-2237, 10'sd384}},
{{11'sd926, 12'sd-1636, 10'sd414}, {10'sd395, 12'sd-1773, 13'sd-2272}, {12'sd-1123, 10'sd-509, 12'sd1729}},
{{13'sd-2171, 13'sd-2579, 12'sd-1516}, {10'sd-467, 12'sd-1202, 12'sd1989}, {12'sd-1092, 12'sd1212, 8'sd108}},
{{11'sd-715, 11'sd-656, 13'sd2724}, {13'sd-2735, 12'sd1496, 12'sd-1344}, {13'sd-2158, 12'sd1194, 12'sd1591}},
{{13'sd2626, 10'sd332, 11'sd-560}, {11'sd801, 12'sd1926, 11'sd-736}, {9'sd-178, 11'sd-616, 13'sd-2880}},
{{12'sd-1341, 10'sd502, 13'sd2178}, {13'sd-2260, 13'sd-2514, 10'sd345}, {13'sd-2103, 13'sd2140, 9'sd200}},
{{12'sd-1120, 12'sd-1634, 8'sd121}, {11'sd859, 12'sd-1558, 11'sd-934}, {10'sd477, 9'sd-174, 13'sd-2577}},
{{9'sd187, 12'sd1359, 13'sd-2801}, {9'sd-166, 12'sd1375, 10'sd401}, {12'sd1277, 11'sd-720, 13'sd-2131}},
{{11'sd-619, 12'sd-1244, 14'sd-4357}, {9'sd-207, 12'sd1808, 10'sd394}, {11'sd-910, 10'sd391, 10'sd412}},
{{11'sd525, 9'sd241, 11'sd-977}, {11'sd-685, 12'sd1192, 13'sd2315}, {13'sd-2182, 13'sd-2677, 13'sd-2501}},
{{9'sd-173, 11'sd748, 5'sd10}, {7'sd-42, 8'sd-79, 13'sd-2709}, {11'sd734, 12'sd1440, 12'sd1228}},
{{12'sd1839, 11'sd838, 12'sd1283}, {13'sd-2300, 13'sd2170, 10'sd-328}, {12'sd1271, 11'sd527, 12'sd1639}},
{{14'sd4207, 11'sd833, 8'sd-108}, {11'sd-838, 12'sd1119, 13'sd-2406}, {13'sd2081, 11'sd-711, 11'sd-904}},
{{11'sd-853, 12'sd-1824, 12'sd-1490}, {11'sd-604, 11'sd678, 12'sd1984}, {12'sd1842, 12'sd-1631, 11'sd-779}},
{{10'sd-267, 12'sd1303, 12'sd1204}, {12'sd2035, 12'sd1324, 10'sd-466}, {11'sd854, 13'sd2363, 12'sd-1777}},
{{13'sd3493, 13'sd3184, 13'sd2048}, {13'sd-2427, 10'sd387, 8'sd106}, {11'sd561, 10'sd-390, 13'sd2439}},
{{12'sd-2026, 12'sd-1656, 13'sd-2809}, {12'sd-1742, 11'sd814, 13'sd-2408}, {13'sd-3451, 12'sd-1539, 9'sd-135}},
{{13'sd-2899, 9'sd-138, 14'sd-5310}, {13'sd-2582, 12'sd1249, 13'sd-2597}, {5'sd10, 13'sd3375, 6'sd-25}},
{{11'sd804, 11'sd782, 10'sd485}, {10'sd-435, 13'sd2617, 12'sd1696}, {13'sd-3736, 12'sd1575, 11'sd-1001}},
{{12'sd-1026, 12'sd-1402, 12'sd-1658}, {12'sd-1312, 11'sd-541, 13'sd-2785}, {10'sd288, 11'sd-886, 12'sd1729}},
{{11'sd807, 12'sd-1073, 12'sd1642}, {11'sd-550, 12'sd-1178, 9'sd-242}, {10'sd285, 13'sd-2589, 11'sd-522}},
{{12'sd1387, 12'sd-1436, 10'sd440}, {12'sd1291, 12'sd1611, 12'sd-1405}, {13'sd-2999, 11'sd872, 11'sd-963}},
{{13'sd-2502, 13'sd-2375, 12'sd1144}, {12'sd1353, 12'sd1238, 10'sd-395}, {12'sd1920, 13'sd-2890, 13'sd-2648}},
{{12'sd-1112, 13'sd-2414, 6'sd-29}, {12'sd-1956, 13'sd-2556, 12'sd1542}, {13'sd2841, 12'sd-1574, 12'sd1799}},
{{13'sd2820, 12'sd-1753, 13'sd2579}, {12'sd1050, 12'sd-1242, 12'sd1503}, {13'sd-2241, 12'sd-1988, 12'sd-1796}},
{{12'sd-1138, 11'sd-596, 10'sd-324}, {12'sd-1380, 11'sd868, 13'sd-2981}, {12'sd1447, 13'sd-2130, 10'sd-285}},
{{7'sd-54, 7'sd61, 12'sd1718}, {12'sd2023, 13'sd2296, 13'sd3099}, {10'sd-456, 6'sd-17, 9'sd-252}},
{{12'sd1926, 13'sd2084, 13'sd3746}, {12'sd-1061, 10'sd-297, 13'sd3158}, {12'sd1572, 9'sd247, 13'sd4001}},
{{12'sd1755, 13'sd2222, 12'sd-1395}, {8'sd-108, 12'sd1696, 12'sd-1035}, {11'sd-537, 12'sd1429, 12'sd-1745}},
{{13'sd-3521, 12'sd1823, 12'sd-1950}, {11'sd544, 12'sd1558, 10'sd337}, {13'sd-2966, 10'sd299, 11'sd980}},
{{13'sd2750, 9'sd200, 12'sd1558}, {13'sd-2161, 12'sd1628, 12'sd-1682}, {12'sd-1252, 12'sd1966, 13'sd2214}},
{{12'sd1494, 12'sd-1379, 12'sd1035}, {8'sd-100, 12'sd1233, 12'sd1650}, {10'sd-346, 13'sd2536, 12'sd-1269}}},
{
{{10'sd-499, 12'sd-1536, 10'sd-349}, {12'sd-1686, 12'sd1647, 12'sd1202}, {13'sd-2614, 11'sd775, 13'sd2221}},
{{13'sd2099, 13'sd-2635, 12'sd-1832}, {12'sd-1940, 10'sd-482, 12'sd1043}, {13'sd2204, 11'sd-766, 12'sd1914}},
{{13'sd2106, 13'sd2182, 13'sd-2203}, {13'sd-2262, 13'sd2176, 13'sd2266}, {13'sd-2195, 13'sd-2453, 13'sd-2082}},
{{12'sd-1475, 10'sd-330, 13'sd2533}, {10'sd-433, 11'sd-586, 10'sd-362}, {12'sd1236, 12'sd1876, 13'sd-2244}},
{{10'sd297, 11'sd-777, 11'sd891}, {12'sd-1968, 9'sd-141, 12'sd-1299}, {9'sd-199, 13'sd-2304, 12'sd-1521}},
{{12'sd-1979, 13'sd-2600, 10'sd-417}, {12'sd-1485, 12'sd1642, 11'sd-864}, {12'sd1592, 8'sd-116, 13'sd2589}},
{{8'sd92, 13'sd2165, 13'sd-2470}, {10'sd439, 13'sd2097, 12'sd1163}, {13'sd-2218, 11'sd715, 13'sd-3041}},
{{13'sd-2396, 10'sd372, 12'sd1110}, {10'sd491, 11'sd-793, 13'sd2603}, {12'sd1653, 12'sd-1065, 12'sd-1199}},
{{13'sd-3164, 12'sd1953, 7'sd-49}, {12'sd-1628, 12'sd-1413, 8'sd111}, {10'sd357, 10'sd-434, 12'sd-1371}},
{{10'sd291, 12'sd1610, 12'sd-1860}, {13'sd-2372, 10'sd-492, 10'sd403}, {10'sd-384, 13'sd-2374, 11'sd-933}},
{{12'sd1839, 9'sd254, 13'sd2901}, {11'sd666, 12'sd-1147, 12'sd-1135}, {11'sd-818, 13'sd2652, 11'sd-540}},
{{12'sd-1842, 12'sd-1916, 9'sd-207}, {12'sd-1295, 11'sd968, 12'sd1274}, {12'sd-1348, 12'sd1500, 12'sd-1511}},
{{11'sd-599, 12'sd-1838, 10'sd420}, {13'sd2920, 5'sd-14, 11'sd685}, {12'sd-1994, 12'sd-1454, 13'sd-2790}},
{{13'sd2371, 13'sd2655, 13'sd-2640}, {10'sd-324, 13'sd-2503, 11'sd606}, {8'sd-119, 13'sd2233, 13'sd-2912}},
{{9'sd-158, 12'sd1249, 11'sd944}, {12'sd1029, 8'sd125, 11'sd863}, {12'sd-1585, 11'sd-744, 12'sd-1755}},
{{10'sd481, 9'sd-129, 12'sd2001}, {12'sd1175, 12'sd1878, 13'sd2705}, {10'sd263, 11'sd-788, 10'sd257}},
{{11'sd-615, 6'sd-16, 12'sd-1307}, {8'sd-125, 12'sd1479, 11'sd-902}, {13'sd-2234, 12'sd1240, 12'sd-1652}},
{{13'sd-2311, 12'sd-1808, 13'sd-2725}, {6'sd-29, 13'sd3773, 13'sd2733}, {12'sd-1312, 13'sd2259, 12'sd1982}},
{{13'sd2846, 13'sd2773, 11'sd880}, {12'sd-1196, 12'sd1538, 13'sd2451}, {10'sd-488, 10'sd330, 11'sd644}},
{{12'sd1275, 9'sd-179, 12'sd-1584}, {13'sd2340, 13'sd2491, 12'sd-1067}, {11'sd-525, 11'sd955, 11'sd686}},
{{12'sd-1621, 12'sd1494, 11'sd-839}, {9'sd-254, 10'sd495, 13'sd-2318}, {13'sd-3120, 10'sd324, 12'sd1688}},
{{9'sd251, 12'sd-1320, 12'sd1406}, {13'sd2679, 13'sd-2370, 12'sd-1208}, {13'sd-2767, 11'sd-925, 12'sd-2042}},
{{12'sd-1748, 13'sd-2355, 13'sd2399}, {10'sd393, 12'sd-1888, 11'sd792}, {11'sd-725, 11'sd-543, 13'sd-2389}},
{{12'sd-1571, 12'sd-1029, 12'sd1825}, {11'sd-971, 11'sd-696, 13'sd2413}, {12'sd-1334, 10'sd-387, 10'sd-271}},
{{12'sd-1530, 12'sd1899, 13'sd2622}, {13'sd2408, 10'sd-401, 10'sd-460}, {11'sd-970, 13'sd2261, 11'sd-841}},
{{11'sd-978, 12'sd-1066, 10'sd-447}, {12'sd1944, 13'sd2821, 12'sd1676}, {10'sd-263, 12'sd-1505, 8'sd106}},
{{11'sd-516, 11'sd517, 7'sd57}, {13'sd-2780, 11'sd-587, 13'sd-2539}, {11'sd-970, 12'sd-1753, 12'sd-1612}},
{{12'sd1741, 12'sd1208, 7'sd-52}, {8'sd-123, 12'sd1893, 11'sd-544}, {11'sd-537, 13'sd-2318, 12'sd-2043}},
{{11'sd797, 12'sd1244, 12'sd-1301}, {12'sd1595, 12'sd-1946, 8'sd-126}, {13'sd2127, 12'sd-1903, 11'sd713}},
{{12'sd1669, 13'sd2474, 12'sd-1941}, {11'sd885, 12'sd-1145, 13'sd-2637}, {12'sd-1797, 12'sd1416, 13'sd2738}},
{{10'sd-385, 12'sd-1453, 12'sd1638}, {12'sd-2039, 11'sd-738, 4'sd7}, {12'sd1275, 12'sd-1650, 12'sd1784}},
{{13'sd-2517, 12'sd-1979, 8'sd109}, {13'sd-3158, 11'sd-538, 11'sd878}, {10'sd-489, 12'sd-1786, 11'sd671}},
{{12'sd-1684, 11'sd913, 12'sd-1084}, {12'sd-1432, 11'sd893, 13'sd-2699}, {13'sd2362, 13'sd2432, 13'sd-2182}},
{{12'sd-1410, 12'sd-1192, 14'sd4133}, {12'sd-1541, 13'sd-2236, 13'sd2692}, {10'sd259, 12'sd1741, 13'sd2310}},
{{13'sd2454, 10'sd304, 12'sd1677}, {12'sd-1371, 13'sd-2172, 13'sd2120}, {13'sd-2642, 11'sd-696, 12'sd1501}},
{{12'sd1969, 13'sd2383, 13'sd2762}, {11'sd1009, 8'sd-86, 12'sd-1209}, {12'sd-1856, 3'sd2, 13'sd2630}},
{{11'sd-691, 13'sd-2788, 10'sd-488}, {13'sd-2945, 10'sd400, 13'sd-2351}, {12'sd1956, 12'sd-1603, 12'sd1269}},
{{12'sd1750, 13'sd2297, 12'sd-1943}, {12'sd1541, 11'sd972, 13'sd2592}, {11'sd-599, 9'sd168, 11'sd-551}},
{{11'sd604, 11'sd-956, 13'sd-2330}, {12'sd1441, 11'sd-705, 10'sd426}, {13'sd2680, 12'sd-1424, 12'sd-1399}},
{{11'sd543, 13'sd-2063, 13'sd2246}, {12'sd-1762, 13'sd2175, 12'sd-1654}, {12'sd1269, 13'sd2463, 12'sd2015}},
{{12'sd-1702, 11'sd-755, 11'sd-822}, {13'sd-3423, 8'sd114, 12'sd1662}, {13'sd-3637, 10'sd303, 10'sd-493}},
{{11'sd-858, 12'sd1478, 13'sd-2812}, {11'sd-861, 8'sd-104, 11'sd915}, {12'sd1589, 12'sd-1514, 12'sd1579}},
{{13'sd-2455, 11'sd-591, 12'sd-1871}, {10'sd262, 13'sd-2345, 12'sd-1625}, {9'sd-206, 12'sd-1694, 13'sd-2847}},
{{12'sd-1298, 11'sd-873, 13'sd2415}, {13'sd2243, 11'sd-950, 13'sd2459}, {9'sd225, 10'sd283, 13'sd2577}},
{{13'sd2119, 8'sd-93, 13'sd2483}, {12'sd-1417, 11'sd763, 12'sd-1148}, {11'sd831, 12'sd1257, 13'sd-2262}},
{{10'sd-469, 12'sd1410, 12'sd-1987}, {9'sd-233, 9'sd210, 9'sd-169}, {12'sd-1471, 11'sd-796, 9'sd-227}},
{{12'sd1902, 12'sd1119, 12'sd1795}, {12'sd-2008, 12'sd1767, 12'sd-1673}, {12'sd1702, 13'sd2855, 12'sd-1513}},
{{11'sd599, 11'sd-654, 11'sd-957}, {8'sd-64, 13'sd-2750, 9'sd229}, {13'sd-2094, 11'sd-993, 13'sd-2622}},
{{12'sd1508, 12'sd-1219, 9'sd-142}, {12'sd-1716, 12'sd1397, 11'sd-933}, {11'sd-1009, 12'sd-1570, 12'sd1417}},
{{8'sd88, 12'sd1063, 9'sd-252}, {11'sd-885, 11'sd-779, 12'sd1268}, {13'sd-2251, 10'sd489, 13'sd2078}},
{{10'sd358, 13'sd2270, 11'sd-855}, {12'sd-1947, 9'sd-221, 12'sd1106}, {12'sd1056, 12'sd1611, 5'sd8}},
{{12'sd-1133, 10'sd374, 12'sd1367}, {12'sd-1065, 13'sd-2576, 11'sd-740}, {12'sd1237, 12'sd-1973, 12'sd-1574}},
{{12'sd1538, 12'sd1731, 13'sd2309}, {12'sd1535, 12'sd1993, 11'sd670}, {13'sd2979, 12'sd1936, 7'sd44}},
{{13'sd2286, 13'sd-2101, 1'sd0}, {9'sd218, 12'sd-1431, 12'sd-2026}, {13'sd-2888, 12'sd1724, 12'sd-1245}},
{{12'sd1153, 12'sd1803, 13'sd-2203}, {12'sd1565, 12'sd-1651, 13'sd-2657}, {12'sd-1142, 12'sd2009, 13'sd-2712}},
{{11'sd682, 13'sd2173, 12'sd1444}, {12'sd-1070, 12'sd1414, 12'sd1526}, {12'sd-1464, 12'sd1484, 13'sd-2427}},
{{12'sd-1370, 11'sd-844, 13'sd-2326}, {9'sd249, 10'sd483, 13'sd2680}, {13'sd-2050, 11'sd-820, 13'sd2060}},
{{1'sd0, 13'sd2156, 12'sd1972}, {13'sd2765, 11'sd700, 12'sd1695}, {13'sd2887, 13'sd2319, 11'sd522}},
{{12'sd1038, 12'sd-1051, 10'sd270}, {12'sd1886, 12'sd1117, 12'sd-1811}, {10'sd-361, 12'sd-1671, 10'sd459}},
{{13'sd2586, 13'sd-2192, 12'sd1659}, {11'sd-592, 13'sd2394, 12'sd-1917}, {9'sd250, 10'sd-430, 12'sd1136}},
{{7'sd59, 9'sd-198, 12'sd1911}, {13'sd-2934, 13'sd-2333, 13'sd2167}, {12'sd-1842, 13'sd2631, 12'sd-1350}},
{{12'sd1638, 13'sd2284, 11'sd-999}, {12'sd1545, 13'sd2110, 11'sd663}, {12'sd1791, 12'sd1265, 11'sd-723}},
{{12'sd1194, 12'sd1331, 11'sd-726}, {13'sd2253, 10'sd-354, 11'sd-626}, {9'sd-183, 13'sd2528, 9'sd204}},
{{12'sd-1187, 11'sd960, 10'sd424}, {12'sd-1502, 13'sd-2506, 5'sd15}, {10'sd-300, 12'sd-1176, 6'sd-16}}},
{
{{10'sd341, 9'sd-159, 12'sd-1178}, {12'sd1614, 11'sd685, 11'sd-881}, {12'sd2029, 10'sd366, 11'sd931}},
{{12'sd1855, 10'sd-400, 10'sd-345}, {13'sd-2278, 12'sd-2045, 12'sd1098}, {13'sd-2634, 12'sd1723, 11'sd559}},
{{11'sd552, 12'sd-1780, 12'sd1319}, {12'sd-1931, 9'sd-137, 13'sd2248}, {12'sd-1559, 13'sd-2098, 11'sd679}},
{{10'sd-401, 12'sd-1178, 13'sd2071}, {12'sd-1382, 11'sd-860, 12'sd1072}, {8'sd-104, 13'sd2249, 12'sd-1103}},
{{12'sd-1950, 13'sd-2713, 7'sd-56}, {7'sd60, 11'sd705, 13'sd2368}, {12'sd-1235, 11'sd953, 11'sd1011}},
{{10'sd440, 11'sd525, 13'sd-2235}, {12'sd-1993, 3'sd3, 12'sd-1255}, {12'sd-1199, 12'sd1980, 12'sd-1065}},
{{9'sd-183, 4'sd4, 12'sd1215}, {12'sd1631, 13'sd3003, 11'sd814}, {13'sd2229, 8'sd82, 12'sd2007}},
{{13'sd2356, 8'sd70, 13'sd3402}, {12'sd1850, 11'sd-886, 13'sd-2698}, {2'sd1, 13'sd-2657, 11'sd555}},
{{12'sd-2031, 13'sd3242, 13'sd2766}, {13'sd2647, 13'sd2324, 12'sd1541}, {11'sd-671, 12'sd1341, 12'sd-1062}},
{{12'sd-1846, 13'sd2290, 12'sd1608}, {11'sd-1017, 12'sd1409, 11'sd635}, {8'sd-82, 13'sd-2349, 4'sd7}},
{{12'sd1122, 11'sd-517, 12'sd1776}, {11'sd782, 11'sd833, 12'sd1127}, {12'sd-1927, 12'sd1438, 12'sd1442}},
{{12'sd1383, 12'sd-1445, 11'sd-979}, {9'sd-234, 13'sd-2170, 11'sd635}, {12'sd-1409, 13'sd-2851, 8'sd-87}},
{{9'sd206, 12'sd1219, 13'sd2514}, {13'sd2571, 11'sd865, 12'sd1986}, {12'sd-1108, 12'sd1748, 13'sd2654}},
{{12'sd1383, 12'sd-1582, 11'sd-866}, {10'sd264, 8'sd102, 13'sd-2053}, {13'sd-2095, 13'sd-2476, 13'sd2092}},
{{13'sd2600, 11'sd675, 12'sd-1560}, {10'sd285, 12'sd-1174, 12'sd-1440}, {8'sd-64, 13'sd-2418, 12'sd-1823}},
{{12'sd-1064, 13'sd2459, 12'sd-1590}, {8'sd67, 13'sd-2644, 10'sd-336}, {12'sd1111, 12'sd-1539, 12'sd1495}},
{{10'sd463, 12'sd1877, 13'sd2137}, {12'sd1927, 12'sd1616, 13'sd-2416}, {9'sd-199, 13'sd-2524, 13'sd2283}},
{{13'sd-2223, 12'sd-1293, 13'sd-3003}, {13'sd2193, 9'sd197, 9'sd-205}, {13'sd2512, 11'sd-987, 13'sd3796}},
{{13'sd2715, 12'sd1041, 12'sd-1501}, {9'sd202, 10'sd-422, 12'sd-1242}, {12'sd1219, 12'sd-1460, 12'sd-1887}},
{{13'sd2327, 12'sd-1282, 13'sd2902}, {12'sd-1771, 13'sd2956, 11'sd918}, {12'sd-1092, 12'sd1887, 11'sd-796}},
{{10'sd-501, 12'sd1744, 12'sd1788}, {13'sd3103, 12'sd-1072, 12'sd1935}, {12'sd-1547, 7'sd60, 11'sd795}},
{{12'sd-1612, 12'sd-1116, 12'sd1703}, {13'sd-2972, 12'sd-1491, 12'sd-1445}, {13'sd-2068, 13'sd2288, 12'sd1686}},
{{11'sd1021, 13'sd2587, 12'sd-1677}, {8'sd-106, 13'sd-2121, 11'sd-872}, {13'sd2469, 12'sd1473, 12'sd1682}},
{{11'sd730, 12'sd1188, 5'sd-12}, {12'sd-1991, 13'sd-2525, 13'sd-2127}, {11'sd772, 12'sd-1722, 11'sd984}},
{{9'sd140, 10'sd266, 12'sd1374}, {12'sd1771, 13'sd2919, 12'sd-1297}, {13'sd2508, 12'sd1941, 11'sd554}},
{{10'sd-393, 13'sd2315, 8'sd-79}, {11'sd-970, 13'sd2084, 12'sd1764}, {10'sd-358, 11'sd-537, 12'sd2020}},
{{12'sd1168, 11'sd-837, 12'sd1232}, {13'sd-2952, 11'sd-891, 12'sd1518}, {10'sd-475, 12'sd-1384, 13'sd-2404}},
{{11'sd-645, 11'sd-582, 11'sd773}, {12'sd-1111, 13'sd3141, 10'sd326}, {13'sd2517, 13'sd-2278, 11'sd-519}},
{{13'sd2116, 12'sd1191, 8'sd-97}, {10'sd-370, 13'sd2370, 13'sd2185}, {12'sd1919, 13'sd2262, 13'sd-2173}},
{{9'sd-217, 9'sd233, 13'sd2785}, {12'sd1283, 12'sd-1644, 11'sd738}, {13'sd-2310, 12'sd-1284, 13'sd-2517}},
{{12'sd-1966, 13'sd-3223, 11'sd-547}, {11'sd-655, 11'sd-966, 11'sd-972}, {12'sd1214, 10'sd-317, 12'sd1400}},
{{12'sd-1235, 11'sd-770, 11'sd-1013}, {12'sd-1217, 13'sd-2714, 12'sd-1269}, {13'sd-2705, 10'sd343, 12'sd1747}},
{{12'sd-1660, 10'sd-347, 13'sd-2658}, {11'sd-965, 12'sd1151, 12'sd1318}, {9'sd-221, 10'sd-422, 12'sd-1541}},
{{11'sd842, 12'sd-1372, 12'sd1489}, {12'sd-1966, 11'sd-881, 10'sd442}, {11'sd-992, 12'sd1212, 11'sd-570}},
{{13'sd-2379, 12'sd-2010, 13'sd2397}, {13'sd2506, 10'sd-380, 10'sd-423}, {13'sd-2148, 12'sd-1869, 9'sd-226}},
{{10'sd-323, 12'sd-1427, 12'sd-1594}, {11'sd-666, 12'sd-1841, 12'sd1445}, {13'sd2298, 12'sd1088, 12'sd1042}},
{{10'sd-283, 11'sd-931, 8'sd-107}, {10'sd413, 13'sd-2518, 12'sd1165}, {13'sd-2177, 11'sd644, 12'sd1162}},
{{12'sd-1768, 12'sd-1404, 13'sd2516}, {11'sd-931, 11'sd861, 12'sd1131}, {11'sd905, 12'sd-1308, 8'sd-119}},
{{12'sd-1430, 10'sd-411, 10'sd-470}, {11'sd865, 13'sd-2455, 12'sd-1256}, {10'sd339, 12'sd-1562, 13'sd3059}},
{{13'sd-2324, 12'sd1033, 13'sd2205}, {13'sd-3034, 11'sd642, 12'sd-1240}, {11'sd984, 11'sd-932, 12'sd-1363}},
{{12'sd-1481, 11'sd-741, 10'sd-421}, {11'sd-718, 10'sd302, 9'sd-246}, {13'sd-2660, 12'sd1815, 9'sd-188}},
{{9'sd-148, 12'sd-1506, 11'sd629}, {12'sd-1319, 12'sd1390, 13'sd-2142}, {11'sd-955, 9'sd-169, 12'sd-1141}},
{{13'sd2642, 11'sd-571, 13'sd-3457}, {13'sd-2411, 10'sd-453, 12'sd1718}, {11'sd848, 12'sd1187, 13'sd-2669}},
{{11'sd-610, 12'sd-1557, 11'sd-930}, {12'sd-1381, 11'sd-545, 12'sd1060}, {13'sd2146, 12'sd2000, 13'sd2284}},
{{13'sd2575, 12'sd1245, 11'sd-725}, {11'sd522, 12'sd-1221, 12'sd-1788}, {13'sd-2368, 11'sd-728, 12'sd-1132}},
{{12'sd1213, 12'sd1928, 12'sd1775}, {12'sd1054, 13'sd2342, 11'sd641}, {11'sd899, 11'sd754, 13'sd2339}},
{{12'sd-1854, 12'sd1026, 12'sd-1374}, {12'sd1576, 12'sd-1451, 12'sd-1860}, {12'sd-1358, 9'sd-175, 11'sd719}},
{{12'sd1230, 9'sd198, 12'sd1034}, {11'sd-982, 11'sd-787, 9'sd-231}, {11'sd546, 5'sd15, 13'sd-2738}},
{{13'sd-2460, 12'sd2031, 13'sd2243}, {5'sd8, 13'sd2156, 13'sd2634}, {13'sd-2265, 13'sd-2193, 12'sd1261}},
{{8'sd118, 10'sd396, 12'sd-1380}, {13'sd2572, 9'sd-186, 8'sd-118}, {11'sd-566, 9'sd179, 11'sd-790}},
{{11'sd-610, 13'sd2199, 13'sd-2255}, {12'sd1357, 12'sd-1720, 13'sd-2066}, {12'sd-1218, 12'sd-1961, 13'sd2176}},
{{12'sd1657, 11'sd640, 11'sd-599}, {5'sd-14, 10'sd264, 11'sd841}, {12'sd-1212, 9'sd-156, 11'sd-1015}},
{{13'sd2676, 12'sd2035, 8'sd114}, {11'sd-781, 13'sd-2504, 13'sd-2457}, {12'sd1435, 7'sd44, 13'sd-2464}},
{{12'sd1436, 11'sd579, 11'sd-589}, {12'sd-1808, 12'sd1638, 13'sd-2168}, {13'sd3048, 4'sd-4, 12'sd1944}},
{{10'sd309, 12'sd1372, 12'sd-1615}, {10'sd279, 12'sd1843, 10'sd-466}, {12'sd-1638, 13'sd3065, 11'sd-679}},
{{11'sd-515, 11'sd777, 12'sd-1212}, {12'sd-2001, 8'sd100, 12'sd-1279}, {12'sd1210, 13'sd2533, 12'sd1772}},
{{13'sd2370, 12'sd1161, 12'sd1699}, {12'sd-1829, 9'sd133, 13'sd-2514}, {13'sd-3205, 12'sd1454, 13'sd2683}},
{{11'sd-756, 12'sd1604, 8'sd96}, {13'sd3343, 11'sd760, 12'sd-1435}, {11'sd738, 13'sd2635, 11'sd-982}},
{{12'sd1760, 9'sd-230, 12'sd-1140}, {11'sd-808, 9'sd160, 11'sd-595}, {13'sd-3027, 11'sd945, 13'sd2503}},
{{12'sd-1049, 13'sd2962, 7'sd32}, {11'sd-859, 13'sd2270, 12'sd1254}, {12'sd-1671, 12'sd-1972, 12'sd1930}},
{{12'sd1868, 10'sd-295, 8'sd-90}, {12'sd-2039, 10'sd-461, 13'sd-2162}, {12'sd1516, 13'sd-2332, 13'sd2489}},
{{12'sd1732, 12'sd-1740, 9'sd174}, {12'sd1104, 11'sd-627, 11'sd969}, {12'sd-1111, 10'sd443, 10'sd485}},
{{13'sd3054, 12'sd1663, 13'sd-2589}, {13'sd-2675, 8'sd-104, 12'sd-1415}, {13'sd2729, 11'sd655, 11'sd-747}},
{{12'sd1909, 12'sd-1401, 12'sd-1384}, {9'sd245, 13'sd-2901, 13'sd-2233}, {13'sd-2511, 10'sd-259, 11'sd-758}}},
{
{{9'sd158, 12'sd-1916, 11'sd1021}, {11'sd-975, 13'sd2131, 12'sd-1241}, {10'sd-309, 12'sd1717, 13'sd2842}},
{{12'sd1093, 9'sd-218, 9'sd215}, {5'sd-10, 13'sd-2706, 12'sd1883}, {12'sd1760, 10'sd-371, 13'sd2728}},
{{13'sd2182, 12'sd-1635, 13'sd2290}, {10'sd435, 12'sd-1153, 11'sd-676}, {13'sd-2740, 11'sd590, 13'sd2137}},
{{11'sd-875, 13'sd-2378, 12'sd1279}, {8'sd-84, 13'sd-2727, 10'sd-310}, {13'sd-2223, 10'sd-504, 12'sd1317}},
{{12'sd1164, 12'sd1325, 12'sd-1122}, {12'sd-1193, 12'sd-1205, 12'sd1748}, {9'sd243, 11'sd-809, 13'sd2572}},
{{7'sd48, 11'sd707, 12'sd-1131}, {12'sd-2013, 11'sd-665, 12'sd-1428}, {12'sd-1489, 12'sd-1081, 12'sd2001}},
{{12'sd-1139, 13'sd-2195, 11'sd-732}, {11'sd892, 12'sd1163, 11'sd972}, {13'sd3238, 13'sd3509, 9'sd-219}},
{{12'sd-1173, 10'sd-398, 12'sd1667}, {9'sd211, 12'sd-1277, 12'sd1792}, {12'sd-1965, 12'sd1263, 13'sd2353}},
{{9'sd177, 11'sd550, 11'sd-567}, {9'sd-131, 13'sd-2248, 12'sd-1967}, {13'sd-2454, 13'sd-2688, 12'sd-1125}},
{{12'sd-1221, 11'sd950, 10'sd502}, {10'sd497, 12'sd1581, 10'sd-286}, {12'sd1821, 10'sd-302, 12'sd1239}},
{{12'sd1699, 12'sd-1824, 13'sd-2268}, {12'sd-1228, 11'sd921, 11'sd621}, {11'sd-547, 13'sd-2471, 13'sd2308}},
{{11'sd908, 11'sd971, 12'sd-1351}, {12'sd-1961, 12'sd1705, 12'sd1294}, {12'sd-1753, 9'sd-243, 13'sd-2572}},
{{10'sd444, 12'sd-1382, 12'sd-1816}, {12'sd1973, 12'sd-1343, 13'sd-2077}, {10'sd292, 11'sd-932, 13'sd2472}},
{{10'sd-279, 11'sd-745, 10'sd-501}, {11'sd-788, 11'sd-744, 12'sd1712}, {12'sd-1097, 13'sd2283, 12'sd-1248}},
{{11'sd-889, 12'sd1391, 13'sd-2186}, {12'sd-1717, 11'sd-928, 12'sd1311}, {13'sd-2997, 12'sd-1345, 13'sd-3409}},
{{13'sd-2087, 10'sd314, 12'sd-1799}, {7'sd-36, 10'sd-259, 13'sd2423}, {12'sd1287, 13'sd-2235, 12'sd-1498}},
{{13'sd2233, 13'sd3206, 12'sd-1339}, {13'sd2465, 13'sd3022, 11'sd-516}, {10'sd-474, 10'sd-394, 11'sd-820}},
{{13'sd3333, 11'sd-881, 11'sd-893}, {13'sd2211, 12'sd-1160, 13'sd-3022}, {13'sd3097, 11'sd609, 11'sd655}},
{{12'sd1501, 13'sd-2104, 11'sd-979}, {12'sd-1944, 8'sd83, 12'sd1387}, {9'sd186, 13'sd-2055, 6'sd23}},
{{11'sd-609, 11'sd-705, 10'sd-444}, {10'sd287, 12'sd-1447, 10'sd347}, {12'sd-1959, 11'sd1011, 10'sd-467}},
{{13'sd3340, 4'sd-4, 12'sd1750}, {12'sd1148, 10'sd432, 13'sd3003}, {12'sd1322, 12'sd1651, 12'sd1190}},
{{10'sd494, 12'sd-1626, 12'sd-1289}, {12'sd-1866, 10'sd393, 12'sd1247}, {9'sd-145, 11'sd921, 11'sd711}},
{{12'sd2033, 12'sd-1775, 12'sd-1809}, {7'sd50, 11'sd-562, 11'sd-793}, {13'sd-2795, 13'sd-2757, 13'sd-2842}},
{{13'sd2053, 13'sd2726, 12'sd1595}, {12'sd1470, 12'sd-1563, 10'sd443}, {11'sd-698, 13'sd2274, 12'sd-1854}},
{{9'sd178, 12'sd1712, 12'sd1750}, {12'sd1808, 13'sd-2609, 12'sd-1599}, {11'sd878, 13'sd-2587, 12'sd1296}},
{{13'sd-2660, 12'sd-1745, 13'sd-2109}, {12'sd-1997, 10'sd353, 11'sd-864}, {7'sd-32, 13'sd-2585, 12'sd1029}},
{{10'sd-418, 12'sd1545, 13'sd2890}, {6'sd-28, 12'sd1377, 12'sd-1431}, {13'sd2772, 12'sd2034, 10'sd424}},
{{11'sd642, 12'sd-1068, 12'sd1575}, {12'sd-1677, 12'sd-1914, 11'sd710}, {12'sd2000, 12'sd1198, 12'sd-1229}},
{{10'sd-467, 12'sd1256, 12'sd-1971}, {8'sd-81, 13'sd2407, 12'sd-1456}, {9'sd-146, 12'sd1982, 12'sd1675}},
{{10'sd-371, 12'sd-1309, 13'sd2677}, {10'sd459, 13'sd-2099, 13'sd-2176}, {11'sd749, 12'sd1318, 9'sd-233}},
{{13'sd2975, 12'sd-1996, 10'sd453}, {11'sd860, 11'sd637, 11'sd-819}, {14'sd5204, 13'sd3611, 7'sd36}},
{{12'sd-1161, 13'sd3013, 12'sd1490}, {13'sd2506, 12'sd1744, 13'sd2144}, {13'sd2618, 12'sd1846, 13'sd-2436}},
{{8'sd80, 12'sd-1568, 11'sd947}, {12'sd1570, 13'sd-2343, 10'sd325}, {9'sd-232, 9'sd-236, 12'sd-1237}},
{{12'sd1064, 13'sd-2305, 13'sd-2459}, {12'sd1884, 12'sd-1844, 12'sd1463}, {12'sd1709, 12'sd-1494, 13'sd-3269}},
{{12'sd1161, 12'sd1227, 12'sd-1806}, {11'sd-732, 12'sd-1091, 13'sd-2113}, {12'sd1339, 13'sd2687, 13'sd2470}},
{{12'sd-1984, 12'sd1188, 13'sd-2229}, {13'sd-2733, 13'sd-2874, 10'sd-272}, {11'sd682, 12'sd1187, 12'sd-1031}},
{{12'sd1395, 12'sd-1535, 12'sd-1447}, {11'sd681, 10'sd-492, 10'sd-505}, {13'sd2214, 11'sd948, 12'sd-1863}},
{{13'sd-2219, 12'sd1546, 12'sd-1670}, {12'sd-1641, 13'sd-2805, 13'sd-2460}, {11'sd689, 12'sd1823, 12'sd-1990}},
{{12'sd1278, 12'sd1591, 11'sd584}, {13'sd-2442, 10'sd432, 12'sd1363}, {12'sd1300, 13'sd-2524, 11'sd517}},
{{11'sd-805, 13'sd2641, 11'sd928}, {12'sd1334, 13'sd-2612, 11'sd538}, {11'sd891, 12'sd-1619, 12'sd-1382}},
{{12'sd-1227, 9'sd177, 8'sd-117}, {11'sd885, 8'sd-116, 4'sd5}, {12'sd-1143, 12'sd1090, 11'sd897}},
{{13'sd-2405, 12'sd1799, 10'sd325}, {11'sd599, 12'sd-1052, 11'sd824}, {10'sd405, 10'sd-355, 8'sd64}},
{{13'sd-2279, 11'sd-949, 8'sd84}, {12'sd-1523, 11'sd-914, 13'sd-2070}, {13'sd-2097, 12'sd-1467, 11'sd-793}},
{{11'sd-899, 11'sd940, 12'sd-1423}, {12'sd-1269, 11'sd-797, 11'sd-682}, {12'sd-1050, 13'sd-2475, 8'sd-101}},
{{12'sd-1072, 12'sd-1636, 12'sd-1216}, {9'sd168, 12'sd1862, 13'sd2872}, {12'sd-1958, 13'sd3201, 12'sd-1079}},
{{13'sd-2194, 12'sd1290, 11'sd956}, {13'sd2137, 9'sd-208, 11'sd-693}, {12'sd1907, 10'sd-378, 11'sd629}},
{{12'sd-1988, 12'sd-1522, 11'sd549}, {13'sd-2428, 12'sd-1135, 13'sd2101}, {12'sd1658, 11'sd762, 12'sd1699}},
{{12'sd-1178, 13'sd2871, 11'sd-1011}, {12'sd1895, 13'sd2255, 13'sd2525}, {7'sd59, 12'sd1083, 12'sd-2031}},
{{9'sd140, 12'sd-1439, 11'sd-561}, {12'sd1320, 12'sd-1919, 11'sd-901}, {13'sd2250, 12'sd1603, 6'sd-19}},
{{13'sd2866, 12'sd-1380, 11'sd1022}, {12'sd1979, 13'sd-2766, 11'sd-533}, {13'sd2126, 13'sd-2243, 11'sd578}},
{{13'sd-3460, 7'sd-63, 13'sd2858}, {13'sd-3225, 11'sd-648, 9'sd-141}, {10'sd329, 11'sd-613, 8'sd98}},
{{12'sd-1037, 13'sd-2847, 11'sd765}, {9'sd214, 10'sd-341, 12'sd-1908}, {11'sd-701, 12'sd1214, 12'sd1836}},
{{12'sd1943, 13'sd2327, 10'sd441}, {10'sd-373, 12'sd-1137, 12'sd1078}, {12'sd-2025, 11'sd637, 9'sd-199}},
{{12'sd-1558, 11'sd-590, 12'sd-1725}, {13'sd3047, 11'sd-749, 12'sd-1246}, {11'sd883, 13'sd-2516, 12'sd-1687}},
{{11'sd783, 10'sd369, 11'sd841}, {7'sd33, 10'sd-263, 13'sd3838}, {12'sd1684, 12'sd-1276, 13'sd2610}},
{{13'sd-2781, 11'sd689, 12'sd-1552}, {12'sd-2032, 12'sd1425, 9'sd-244}, {12'sd1972, 10'sd-349, 13'sd-2283}},
{{7'sd-59, 9'sd204, 13'sd2419}, {12'sd1084, 11'sd701, 7'sd54}, {12'sd-1187, 12'sd1385, 11'sd702}},
{{10'sd414, 11'sd854, 13'sd-2067}, {13'sd-2219, 11'sd-702, 13'sd-2318}, {11'sd-741, 12'sd1913, 11'sd-587}},
{{12'sd1285, 13'sd2339, 12'sd-1603}, {12'sd-1694, 7'sd-43, 13'sd2091}, {12'sd-1057, 12'sd1255, 8'sd118}},
{{13'sd2432, 13'sd-2714, 13'sd2821}, {13'sd-2502, 12'sd-1657, 6'sd-20}, {10'sd477, 11'sd909, 13'sd3115}},
{{13'sd2477, 12'sd1194, 9'sd192}, {13'sd2937, 12'sd1413, 12'sd1226}, {12'sd-1556, 12'sd-1187, 13'sd-2065}},
{{13'sd-2239, 12'sd-1351, 10'sd302}, {13'sd2252, 10'sd335, 12'sd1752}, {13'sd2492, 12'sd1694, 13'sd2134}},
{{13'sd-2333, 13'sd-2529, 9'sd-240}, {13'sd2506, 11'sd-967, 12'sd1245}, {12'sd-1555, 11'sd1011, 12'sd1528}},
{{10'sd481, 7'sd36, 11'sd-721}, {13'sd2175, 11'sd924, 11'sd-808}, {10'sd-285, 12'sd-1547, 11'sd620}}},
{
{{8'sd74, 13'sd2712, 11'sd-772}, {12'sd-1909, 10'sd-356, 9'sd-158}, {13'sd2274, 13'sd-2929, 10'sd-284}},
{{13'sd-2882, 12'sd1636, 12'sd-1315}, {12'sd1350, 12'sd-1805, 11'sd542}, {11'sd666, 11'sd644, 12'sd1733}},
{{13'sd2953, 13'sd2370, 13'sd2969}, {12'sd1876, 11'sd-696, 13'sd-2599}, {13'sd-2933, 12'sd1958, 12'sd-1198}},
{{10'sd305, 11'sd-960, 12'sd1112}, {12'sd1572, 8'sd-112, 13'sd-2055}, {13'sd2159, 11'sd-632, 11'sd689}},
{{10'sd-500, 12'sd2009, 12'sd-1511}, {12'sd1145, 11'sd563, 13'sd2910}, {11'sd672, 11'sd-558, 12'sd1840}},
{{12'sd1407, 11'sd-923, 9'sd-160}, {12'sd-1362, 12'sd-1328, 11'sd-556}, {13'sd-2211, 11'sd977, 11'sd715}},
{{12'sd1408, 12'sd-1985, 12'sd-1775}, {12'sd1641, 12'sd1781, 12'sd-1820}, {12'sd1725, 12'sd1620, 8'sd104}},
{{11'sd623, 13'sd2633, 8'sd125}, {13'sd2553, 13'sd2433, 12'sd1076}, {12'sd-1750, 12'sd-1493, 11'sd575}},
{{12'sd-1842, 12'sd1207, 12'sd1353}, {9'sd214, 9'sd-188, 13'sd-3179}, {10'sd-507, 7'sd-50, 9'sd-214}},
{{12'sd-1352, 12'sd1376, 12'sd1045}, {13'sd2149, 10'sd374, 13'sd2348}, {12'sd1515, 8'sd89, 12'sd-1248}},
{{11'sd-992, 11'sd-723, 13'sd-2301}, {13'sd-2709, 12'sd-1446, 8'sd-111}, {12'sd1074, 10'sd398, 13'sd-2761}},
{{12'sd1175, 12'sd-1914, 13'sd-2508}, {13'sd2346, 10'sd283, 8'sd119}, {11'sd585, 12'sd-2007, 10'sd430}},
{{10'sd-447, 12'sd-1620, 11'sd621}, {11'sd629, 13'sd-3685, 13'sd-2242}, {12'sd1848, 13'sd2287, 11'sd591}},
{{13'sd-2990, 11'sd570, 13'sd2208}, {12'sd1949, 12'sd1256, 12'sd-1554}, {11'sd674, 10'sd329, 13'sd-2845}},
{{11'sd-767, 11'sd558, 13'sd2601}, {6'sd-25, 13'sd2886, 12'sd-1792}, {13'sd-2856, 12'sd1431, 9'sd-240}},
{{12'sd1934, 11'sd642, 12'sd-1464}, {11'sd-851, 12'sd-1591, 8'sd95}, {8'sd-92, 13'sd2559, 10'sd-439}},
{{13'sd-2336, 13'sd-2125, 12'sd1036}, {13'sd2127, 11'sd879, 13'sd2485}, {12'sd1935, 11'sd969, 13'sd2637}},
{{13'sd2299, 11'sd914, 12'sd1783}, {12'sd1281, 12'sd-1813, 13'sd-2177}, {13'sd2856, 13'sd-2705, 12'sd-1547}},
{{11'sd-865, 11'sd-786, 6'sd-29}, {11'sd-1023, 13'sd2500, 12'sd-1764}, {10'sd470, 8'sd-113, 6'sd-17}},
{{13'sd-2308, 13'sd-2843, 13'sd-2716}, {13'sd-2349, 11'sd-519, 13'sd-2751}, {12'sd-1736, 11'sd-696, 12'sd-2042}},
{{10'sd399, 13'sd-2716, 11'sd-713}, {12'sd-1179, 12'sd1523, 11'sd-831}, {12'sd-1384, 10'sd314, 13'sd-2661}},
{{11'sd676, 10'sd-273, 12'sd-1500}, {12'sd-1436, 11'sd-698, 12'sd-1565}, {13'sd-2152, 12'sd1444, 11'sd-740}},
{{12'sd1888, 11'sd-777, 12'sd-2030}, {12'sd1546, 13'sd2135, 10'sd-276}, {12'sd1948, 10'sd340, 12'sd1257}},
{{6'sd18, 12'sd1053, 13'sd-2244}, {12'sd-1756, 13'sd3023, 12'sd-1159}, {11'sd780, 9'sd-175, 11'sd-731}},
{{12'sd1516, 12'sd1240, 13'sd-2152}, {12'sd-1576, 13'sd-2160, 10'sd-315}, {13'sd-2283, 11'sd982, 11'sd-984}},
{{12'sd1303, 9'sd170, 12'sd-1952}, {13'sd-2389, 13'sd-2659, 12'sd-1800}, {12'sd-1945, 13'sd-2705, 12'sd1930}},
{{12'sd1257, 9'sd-141, 12'sd-1866}, {13'sd2796, 13'sd-2299, 13'sd2052}, {12'sd1139, 12'sd-2005, 12'sd-1750}},
{{13'sd-2935, 12'sd1738, 13'sd2739}, {11'sd937, 8'sd69, 12'sd-1099}, {10'sd-321, 6'sd23, 6'sd-30}},
{{13'sd-2181, 13'sd-2735, 13'sd2408}, {11'sd689, 9'sd-206, 12'sd-1122}, {12'sd1221, 11'sd-545, 9'sd-219}},
{{11'sd694, 12'sd-1364, 13'sd2343}, {12'sd1846, 13'sd-2301, 12'sd-1282}, {12'sd-1625, 8'sd-117, 12'sd1891}},
{{11'sd-542, 12'sd1445, 12'sd-1630}, {12'sd-1783, 12'sd-1376, 13'sd2563}, {13'sd3023, 10'sd481, 11'sd-965}},
{{13'sd2760, 12'sd-1765, 9'sd215}, {13'sd2501, 11'sd642, 12'sd1107}, {11'sd590, 12'sd-1211, 13'sd2360}},
{{12'sd1501, 12'sd-1545, 13'sd2324}, {11'sd-809, 12'sd-1261, 13'sd2170}, {7'sd41, 12'sd1345, 9'sd-152}},
{{12'sd1802, 11'sd-536, 9'sd-224}, {12'sd-1533, 13'sd2454, 9'sd-202}, {10'sd-434, 8'sd120, 10'sd356}},
{{12'sd1365, 11'sd574, 12'sd-1707}, {12'sd1064, 11'sd-789, 11'sd722}, {12'sd-1678, 12'sd1329, 12'sd1443}},
{{12'sd-1160, 12'sd-1615, 10'sd295}, {10'sd365, 9'sd-197, 13'sd-2794}, {10'sd-270, 12'sd1753, 13'sd-2293}},
{{11'sd-590, 9'sd140, 13'sd-2373}, {13'sd-2260, 12'sd1353, 13'sd-2707}, {11'sd745, 12'sd1615, 13'sd-3048}},
{{13'sd-2276, 12'sd1202, 11'sd-717}, {12'sd-1556, 11'sd697, 8'sd98}, {9'sd211, 12'sd-1184, 11'sd-619}},
{{12'sd1837, 12'sd-1183, 12'sd1638}, {12'sd-1154, 12'sd-1253, 12'sd1867}, {12'sd-2046, 13'sd-2581, 13'sd2134}},
{{6'sd-17, 11'sd-810, 12'sd1591}, {12'sd-1182, 11'sd-835, 13'sd-2452}, {11'sd614, 11'sd759, 12'sd1711}},
{{13'sd-2212, 12'sd1163, 12'sd-1158}, {13'sd-2216, 12'sd1117, 13'sd-2229}, {13'sd-2835, 11'sd-930, 13'sd-2645}},
{{12'sd1179, 11'sd793, 10'sd448}, {13'sd-2501, 11'sd-780, 12'sd-1119}, {8'sd65, 3'sd-3, 13'sd2338}},
{{10'sd-386, 13'sd2204, 12'sd1626}, {13'sd-3195, 12'sd1859, 12'sd-1207}, {13'sd-2694, 13'sd-2147, 13'sd2526}},
{{9'sd-218, 11'sd964, 12'sd-1835}, {13'sd-3041, 9'sd-173, 12'sd1382}, {12'sd1373, 9'sd-182, 12'sd1659}},
{{12'sd1158, 12'sd-1457, 12'sd1480}, {13'sd-2687, 13'sd2713, 10'sd324}, {13'sd-2557, 11'sd-817, 13'sd2526}},
{{12'sd1284, 12'sd1099, 12'sd-1832}, {9'sd-222, 12'sd-2005, 13'sd-2162}, {13'sd-2821, 10'sd276, 12'sd1896}},
{{12'sd1089, 12'sd-1770, 13'sd-2637}, {13'sd-2196, 12'sd1903, 13'sd2055}, {13'sd-2699, 13'sd-3096, 13'sd-2819}},
{{12'sd1354, 8'sd69, 10'sd511}, {12'sd-1202, 11'sd928, 12'sd1576}, {12'sd1475, 12'sd-1079, 13'sd3305}},
{{13'sd3843, 12'sd-1544, 13'sd-3078}, {12'sd1643, 13'sd2505, 11'sd587}, {13'sd2320, 12'sd1327, 13'sd-2612}},
{{8'sd-76, 12'sd1946, 10'sd-263}, {12'sd1769, 12'sd-1347, 13'sd2559}, {12'sd2009, 11'sd981, 8'sd87}},
{{12'sd-1976, 13'sd2098, 9'sd215}, {11'sd-904, 11'sd-760, 13'sd3703}, {14'sd-4310, 11'sd772, 13'sd2352}},
{{12'sd1921, 12'sd1719, 11'sd-882}, {12'sd1330, 10'sd401, 12'sd1486}, {11'sd-633, 13'sd-2835, 11'sd-946}},
{{11'sd577, 11'sd662, 13'sd-2133}, {13'sd-2452, 12'sd-1040, 10'sd-306}, {13'sd-2171, 12'sd1761, 6'sd21}},
{{12'sd-1133, 12'sd1103, 13'sd2823}, {12'sd-1601, 5'sd14, 11'sd895}, {11'sd-741, 13'sd2182, 10'sd432}},
{{13'sd2559, 13'sd-2068, 13'sd3813}, {13'sd-3220, 12'sd-1819, 9'sd-164}, {13'sd2532, 12'sd-1721, 8'sd-122}},
{{13'sd2173, 13'sd-2382, 13'sd-2512}, {13'sd-2145, 9'sd-132, 12'sd2044}, {13'sd2108, 13'sd-2334, 13'sd2633}},
{{13'sd2302, 12'sd-1234, 7'sd-48}, {10'sd-290, 13'sd-2056, 11'sd-571}, {12'sd1530, 11'sd-599, 12'sd-1642}},
{{12'sd-1860, 13'sd-2112, 10'sd-502}, {11'sd914, 12'sd1178, 10'sd359}, {11'sd832, 12'sd2044, 13'sd2337}},
{{10'sd341, 11'sd654, 13'sd-2210}, {11'sd594, 13'sd-2222, 12'sd1106}, {13'sd-2431, 12'sd-1572, 11'sd-788}},
{{12'sd1291, 10'sd-304, 13'sd3490}, {11'sd-797, 12'sd-1487, 12'sd-1558}, {12'sd-1328, 12'sd-1275, 12'sd-1264}},
{{12'sd-1508, 10'sd-339, 12'sd1236}, {9'sd177, 12'sd1749, 12'sd1877}, {13'sd2487, 11'sd-990, 13'sd-2282}},
{{12'sd-1989, 12'sd-1504, 11'sd622}, {13'sd-2076, 12'sd-1712, 12'sd-1444}, {12'sd1177, 13'sd-2276, 12'sd-1844}},
{{8'sd-105, 10'sd-308, 9'sd132}, {13'sd2373, 12'sd1880, 13'sd2360}, {11'sd-781, 11'sd921, 13'sd2433}},
{{13'sd2602, 12'sd1260, 9'sd134}, {13'sd2606, 11'sd-705, 12'sd1391}, {12'sd-1043, 13'sd-2076, 10'sd-349}}},
{
{{13'sd-2838, 4'sd4, 12'sd-1880}, {12'sd-1886, 13'sd2620, 12'sd-1829}, {13'sd-2819, 11'sd-665, 12'sd1375}},
{{13'sd-2774, 10'sd-490, 13'sd-2055}, {12'sd1219, 11'sd531, 13'sd2202}, {11'sd756, 13'sd-2274, 6'sd21}},
{{11'sd-758, 12'sd-1589, 13'sd-2279}, {12'sd1061, 12'sd-1084, 8'sd-126}, {13'sd-2562, 12'sd1460, 12'sd-1936}},
{{12'sd-1460, 13'sd-2227, 13'sd-3238}, {11'sd680, 13'sd-2473, 12'sd-1827}, {13'sd-2997, 12'sd1911, 10'sd441}},
{{12'sd1611, 12'sd-2019, 13'sd2458}, {12'sd-1480, 12'sd1720, 12'sd-1574}, {10'sd471, 12'sd-1701, 11'sd724}},
{{12'sd-1751, 13'sd2199, 13'sd2589}, {10'sd-290, 10'sd-382, 12'sd1206}, {13'sd2570, 12'sd1040, 11'sd919}},
{{13'sd-3059, 11'sd791, 10'sd484}, {11'sd-557, 12'sd-1233, 12'sd-1921}, {9'sd-182, 13'sd2804, 11'sd-983}},
{{12'sd1329, 12'sd-1330, 10'sd451}, {12'sd-1986, 11'sd885, 4'sd6}, {12'sd-1058, 7'sd38, 12'sd1468}},
{{13'sd2994, 13'sd-2787, 11'sd973}, {12'sd1993, 12'sd-1417, 9'sd168}, {12'sd-1920, 12'sd-2028, 10'sd346}},
{{12'sd-1462, 11'sd-770, 13'sd2636}, {12'sd1426, 13'sd2818, 11'sd752}, {13'sd-2571, 13'sd2565, 13'sd2178}},
{{11'sd-1005, 12'sd1418, 8'sd83}, {12'sd-2006, 12'sd-1999, 12'sd1437}, {10'sd458, 12'sd1618, 12'sd-1481}},
{{11'sd-890, 12'sd-1267, 11'sd-903}, {11'sd923, 12'sd-1117, 12'sd-1923}, {12'sd2010, 12'sd1920, 11'sd569}},
{{12'sd-1259, 12'sd-1890, 13'sd-2392}, {11'sd-586, 12'sd1867, 13'sd-2303}, {13'sd2051, 12'sd-1404, 13'sd2116}},
{{13'sd-2716, 13'sd-2155, 12'sd-1985}, {12'sd-1078, 13'sd-2477, 10'sd-414}, {12'sd1273, 11'sd978, 11'sd606}},
{{13'sd2144, 11'sd778, 13'sd2169}, {11'sd-529, 13'sd-2053, 13'sd2340}, {13'sd-2792, 13'sd2171, 9'sd202}},
{{12'sd1133, 11'sd633, 13'sd-2437}, {12'sd-1343, 12'sd1197, 12'sd1763}, {13'sd2090, 12'sd1936, 12'sd-1879}},
{{11'sd660, 7'sd-35, 10'sd286}, {13'sd2390, 9'sd-213, 13'sd-2376}, {12'sd1335, 13'sd-2051, 13'sd2276}},
{{6'sd-20, 13'sd2389, 13'sd-3277}, {12'sd-1419, 12'sd1234, 11'sd-523}, {12'sd-1162, 10'sd-375, 12'sd-1891}},
{{13'sd2322, 13'sd-2521, 9'sd132}, {11'sd546, 13'sd-2075, 10'sd266}, {12'sd1590, 13'sd2753, 12'sd1421}},
{{12'sd-1498, 9'sd-156, 11'sd-742}, {12'sd-1088, 13'sd-3181, 13'sd-2742}, {12'sd-1172, 13'sd-2822, 12'sd-1802}},
{{11'sd-826, 13'sd-2217, 11'sd663}, {12'sd1212, 12'sd1309, 13'sd-2595}, {12'sd-1761, 11'sd-931, 12'sd-1439}},
{{11'sd743, 11'sd-799, 13'sd-2750}, {12'sd1431, 11'sd703, 8'sd-117}, {10'sd395, 13'sd2375, 13'sd-2591}},
{{12'sd-1179, 13'sd-2243, 10'sd-393}, {13'sd2806, 13'sd2070, 12'sd-1358}, {12'sd1316, 12'sd-1446, 12'sd1799}},
{{12'sd-1285, 13'sd3139, 11'sd761}, {11'sd969, 12'sd1493, 12'sd1429}, {12'sd-1882, 13'sd2430, 10'sd460}},
{{11'sd-804, 13'sd2148, 13'sd-2532}, {12'sd-1324, 11'sd685, 13'sd2354}, {12'sd-1429, 12'sd-1052, 11'sd766}},
{{12'sd1060, 9'sd-231, 12'sd1757}, {13'sd-2424, 13'sd2149, 13'sd-2110}, {11'sd717, 10'sd263, 13'sd-2586}},
{{12'sd1159, 13'sd3086, 13'sd2254}, {12'sd1227, 10'sd339, 13'sd2364}, {12'sd-1942, 11'sd-947, 12'sd1955}},
{{13'sd-2555, 10'sd369, 10'sd454}, {9'sd-148, 12'sd1364, 13'sd2419}, {11'sd-933, 12'sd1307, 12'sd1935}},
{{11'sd-964, 13'sd2238, 11'sd-688}, {12'sd1850, 12'sd-1565, 13'sd2118}, {13'sd2126, 13'sd-2099, 13'sd2223}},
{{13'sd2560, 11'sd542, 13'sd2501}, {11'sd947, 13'sd-2075, 13'sd-2458}, {13'sd-2167, 12'sd-1515, 8'sd93}},
{{12'sd-1119, 7'sd53, 8'sd108}, {10'sd302, 12'sd-1873, 11'sd-966}, {14'sd4524, 13'sd3337, 11'sd-516}},
{{11'sd-670, 13'sd-2191, 12'sd1363}, {12'sd1364, 11'sd-737, 12'sd1342}, {12'sd1625, 12'sd-1445, 12'sd1570}},
{{12'sd2000, 12'sd1346, 11'sd838}, {10'sd463, 12'sd-1445, 13'sd-2212}, {7'sd-44, 12'sd1155, 11'sd550}},
{{10'sd-322, 11'sd-766, 10'sd-352}, {12'sd1796, 13'sd2170, 10'sd-323}, {13'sd3133, 12'sd1212, 12'sd1886}},
{{12'sd-1278, 13'sd2226, 13'sd2659}, {13'sd-2543, 10'sd309, 10'sd-266}, {12'sd-1122, 12'sd1481, 13'sd-2187}},
{{13'sd-2837, 11'sd798, 11'sd712}, {9'sd248, 12'sd1683, 13'sd2285}, {7'sd-48, 13'sd-2696, 12'sd-1265}},
{{9'sd-218, 5'sd-13, 12'sd-1847}, {11'sd-941, 11'sd707, 13'sd2381}, {11'sd741, 12'sd-1366, 13'sd2224}},
{{11'sd-931, 12'sd1363, 13'sd-2898}, {12'sd1078, 13'sd-2343, 12'sd1336}, {13'sd2674, 13'sd-2668, 11'sd-677}},
{{12'sd1946, 12'sd-1428, 13'sd-2247}, {12'sd1058, 11'sd-988, 11'sd840}, {9'sd-211, 11'sd816, 10'sd-260}},
{{8'sd-98, 13'sd-2082, 12'sd1398}, {11'sd-585, 13'sd2636, 10'sd511}, {13'sd2348, 10'sd262, 13'sd-2743}},
{{11'sd-615, 7'sd56, 12'sd1793}, {7'sd-35, 13'sd2090, 12'sd1971}, {12'sd-1445, 11'sd-656, 10'sd-352}},
{{12'sd-1172, 12'sd-2044, 13'sd2568}, {12'sd1302, 12'sd-1670, 13'sd3043}, {13'sd2331, 11'sd534, 12'sd1845}},
{{9'sd-196, 11'sd912, 13'sd-2105}, {13'sd-2588, 8'sd87, 13'sd-2075}, {12'sd-1635, 12'sd-1757, 9'sd185}},
{{13'sd-2805, 13'sd-3050, 11'sd705}, {9'sd208, 13'sd-2206, 8'sd-112}, {13'sd-2774, 13'sd-2609, 9'sd-243}},
{{11'sd930, 12'sd1348, 12'sd1233}, {12'sd-2045, 12'sd-1965, 11'sd799}, {13'sd-2717, 11'sd-928, 10'sd-437}},
{{11'sd-952, 10'sd-294, 11'sd714}, {13'sd2177, 12'sd-1677, 13'sd2142}, {13'sd-2553, 13'sd-2958, 12'sd1574}},
{{8'sd-115, 10'sd302, 12'sd-1298}, {12'sd-1382, 12'sd-1998, 13'sd-2097}, {12'sd2022, 9'sd197, 13'sd-2048}},
{{12'sd-1920, 13'sd-2736, 13'sd2501}, {13'sd-2322, 13'sd-2302, 13'sd2729}, {12'sd1275, 13'sd3169, 7'sd-54}},
{{13'sd2909, 11'sd-711, 13'sd-2468}, {13'sd2693, 11'sd-562, 12'sd1364}, {8'sd-66, 13'sd-2430, 10'sd333}},
{{12'sd1680, 12'sd1640, 12'sd1238}, {7'sd38, 6'sd23, 11'sd-891}, {6'sd26, 12'sd-2003, 12'sd-1428}},
{{13'sd-2127, 12'sd1664, 13'sd2221}, {6'sd-23, 13'sd2226, 11'sd851}, {13'sd-3873, 12'sd-1299, 12'sd-1129}},
{{13'sd-2630, 13'sd-2221, 11'sd886}, {9'sd174, 12'sd1565, 12'sd1790}, {12'sd1685, 11'sd740, 12'sd-1409}},
{{12'sd1598, 13'sd-2079, 10'sd291}, {13'sd-2677, 13'sd-2458, 13'sd-2748}, {13'sd2672, 13'sd-2402, 12'sd-1255}},
{{12'sd1575, 12'sd-1874, 13'sd2151}, {13'sd-2243, 10'sd344, 11'sd-842}, {11'sd-999, 12'sd-1722, 9'sd180}},
{{12'sd-1107, 12'sd1357, 9'sd-245}, {11'sd836, 10'sd329, 11'sd800}, {11'sd-839, 10'sd320, 12'sd-1889}},
{{13'sd-2468, 12'sd-1558, 12'sd1438}, {13'sd-2644, 11'sd914, 12'sd1026}, {9'sd-207, 11'sd-904, 11'sd746}},
{{12'sd1322, 10'sd-408, 10'sd305}, {11'sd964, 12'sd1753, 10'sd-455}, {10'sd479, 13'sd2784, 13'sd2551}},
{{11'sd618, 13'sd2738, 11'sd-720}, {10'sd-504, 12'sd-1305, 12'sd1293}, {11'sd-641, 12'sd2005, 11'sd1016}},
{{13'sd-2302, 11'sd-580, 11'sd-879}, {12'sd-2029, 13'sd2865, 12'sd-1103}, {12'sd1426, 13'sd-2048, 13'sd2694}},
{{12'sd1142, 11'sd702, 13'sd2424}, {11'sd-515, 12'sd-1279, 13'sd2618}, {12'sd1286, 12'sd-1672, 11'sd-801}},
{{12'sd1799, 10'sd-467, 12'sd1697}, {11'sd-573, 13'sd3062, 11'sd574}, {12'sd1934, 12'sd1899, 11'sd592}},
{{13'sd-2501, 12'sd1317, 11'sd975}, {11'sd839, 12'sd1220, 12'sd-1290}, {13'sd3016, 9'sd192, 6'sd21}},
{{13'sd-2077, 12'sd1296, 12'sd1870}, {11'sd-606, 12'sd1112, 13'sd2230}, {12'sd-1268, 12'sd1623, 9'sd-252}},
{{13'sd-2100, 12'sd1242, 13'sd-3226}, {12'sd1841, 10'sd-263, 12'sd1695}, {13'sd-2201, 12'sd-1384, 13'sd-2387}}}},
// Weights for conv5_weight
{
{
{{12'sd1699, 11'sd540, 12'sd-1847}, {12'sd-1985, 13'sd2074, 13'sd2618}, {7'sd54, 11'sd-879, 11'sd948}},
{{12'sd1461, 11'sd560, 11'sd562}, {12'sd1422, 13'sd2530, 13'sd2483}, {9'sd191, 10'sd309, 13'sd3630}},
{{12'sd1113, 13'sd2244, 12'sd-1862}, {12'sd1362, 10'sd-365, 13'sd2474}, {13'sd-2182, 12'sd-1153, 9'sd172}},
{{11'sd-823, 11'sd593, 11'sd600}, {12'sd1663, 13'sd2941, 11'sd-609}, {11'sd-903, 12'sd-1414, 11'sd-920}},
{{8'sd105, 7'sd47, 12'sd1180}, {11'sd887, 11'sd-680, 5'sd-12}, {12'sd1909, 12'sd-1527, 11'sd689}},
{{13'sd2248, 11'sd658, 13'sd2115}, {8'sd97, 12'sd-1048, 13'sd2231}, {13'sd2317, 11'sd670, 13'sd2580}},
{{11'sd-859, 12'sd1183, 10'sd297}, {10'sd449, 13'sd2846, 12'sd-1733}, {12'sd-1729, 12'sd-1595, 11'sd-904}},
{{11'sd952, 11'sd998, 13'sd-2792}, {13'sd2061, 13'sd3005, 10'sd511}, {13'sd3358, 12'sd-1410, 12'sd-1781}},
{{13'sd2313, 12'sd-1617, 13'sd2296}, {12'sd-1268, 12'sd-1141, 12'sd-1667}, {11'sd757, 9'sd134, 11'sd608}},
{{12'sd1445, 11'sd768, 9'sd-170}, {9'sd232, 9'sd-206, 12'sd1028}, {12'sd-1752, 11'sd773, 8'sd69}},
{{13'sd-2573, 10'sd-454, 13'sd-2380}, {12'sd-1887, 12'sd-1993, 11'sd1005}, {12'sd-1851, 13'sd-2815, 12'sd-2028}},
{{12'sd-1346, 12'sd1898, 10'sd-482}, {11'sd834, 11'sd816, 11'sd-703}, {11'sd1020, 10'sd293, 11'sd-779}},
{{12'sd1442, 12'sd-1286, 12'sd1787}, {12'sd1183, 9'sd173, 13'sd-2103}, {11'sd-638, 12'sd1342, 12'sd-1717}},
{{13'sd-2999, 12'sd-1681, 9'sd208}, {10'sd-408, 12'sd1106, 11'sd702}, {9'sd-182, 12'sd1943, 10'sd-395}},
{{13'sd-2515, 12'sd-1300, 12'sd1302}, {11'sd-700, 13'sd2619, 13'sd2128}, {13'sd-3803, 12'sd1711, 10'sd266}},
{{11'sd-755, 12'sd-1462, 11'sd852}, {12'sd1854, 12'sd-1625, 8'sd-98}, {11'sd-547, 11'sd-815, 11'sd987}},
{{12'sd-1520, 12'sd-2017, 12'sd1110}, {12'sd1608, 11'sd-988, 11'sd787}, {12'sd-1911, 12'sd1315, 13'sd2188}},
{{12'sd1500, 10'sd-334, 13'sd2918}, {12'sd1129, 12'sd1618, 13'sd2214}, {12'sd1786, 12'sd-1474, 11'sd742}},
{{13'sd-2309, 13'sd2051, 12'sd1443}, {13'sd2907, 12'sd2044, 12'sd1356}, {13'sd2773, 10'sd-314, 10'sd-318}},
{{13'sd-2410, 11'sd554, 11'sd864}, {13'sd2236, 11'sd-542, 13'sd-2430}, {13'sd2261, 12'sd1332, 10'sd-324}},
{{12'sd1049, 13'sd2809, 12'sd1547}, {12'sd2010, 12'sd-1472, 12'sd1429}, {13'sd-2625, 13'sd-2071, 13'sd-2234}},
{{14'sd4153, 12'sd1728, 12'sd-1762}, {11'sd752, 12'sd-1718, 12'sd2031}, {13'sd-2273, 13'sd-2881, 11'sd-705}},
{{9'sd-152, 8'sd-98, 13'sd-2882}, {11'sd818, 12'sd-1655, 13'sd-2612}, {11'sd624, 11'sd957, 11'sd-675}},
{{12'sd1796, 10'sd367, 12'sd1270}, {10'sd-408, 12'sd-1911, 12'sd-1137}, {12'sd1294, 11'sd616, 13'sd-3947}},
{{13'sd-2158, 12'sd1983, 13'sd3235}, {12'sd1172, 13'sd-2613, 12'sd-1514}, {12'sd1271, 10'sd-345, 11'sd-546}},
{{13'sd-2256, 11'sd-516, 13'sd-3050}, {12'sd1765, 12'sd1409, 11'sd967}, {13'sd2998, 12'sd1236, 13'sd-2091}},
{{12'sd1485, 13'sd-2609, 13'sd-2211}, {11'sd838, 13'sd-2492, 9'sd196}, {11'sd-728, 13'sd-2798, 12'sd1973}},
{{12'sd1181, 11'sd561, 12'sd1026}, {13'sd-2144, 10'sd-309, 8'sd100}, {13'sd-3200, 11'sd859, 12'sd1151}},
{{12'sd-2030, 12'sd1269, 7'sd51}, {12'sd-1328, 10'sd503, 12'sd1897}, {11'sd891, 11'sd663, 10'sd-273}},
{{13'sd2964, 12'sd1612, 12'sd-1217}, {13'sd3116, 13'sd2374, 12'sd1638}, {13'sd3023, 13'sd2133, 13'sd2859}},
{{12'sd-1998, 12'sd1248, 13'sd-2755}, {12'sd1963, 12'sd1564, 12'sd1290}, {12'sd-1816, 9'sd-208, 12'sd2025}},
{{10'sd480, 11'sd-904, 11'sd-549}, {12'sd1648, 12'sd1994, 11'sd-879}, {11'sd736, 12'sd-1940, 13'sd-2053}},
{{11'sd797, 12'sd2032, 13'sd2067}, {13'sd-2855, 13'sd2194, 13'sd-2979}, {13'sd2430, 13'sd2422, 12'sd-1656}},
{{12'sd1201, 12'sd1115, 13'sd2426}, {12'sd1168, 12'sd1552, 12'sd1056}, {13'sd-2394, 12'sd-1194, 11'sd-779}},
{{12'sd1271, 12'sd-1991, 13'sd-3553}, {13'sd2167, 12'sd1971, 13'sd-2989}, {14'sd4117, 7'sd58, 13'sd-2055}},
{{11'sd-819, 12'sd2036, 12'sd1222}, {11'sd-793, 10'sd-510, 10'sd415}, {11'sd896, 13'sd2195, 12'sd1244}},
{{12'sd-1206, 10'sd-261, 12'sd1220}, {13'sd2869, 12'sd1375, 12'sd1984}, {13'sd2757, 13'sd3055, 13'sd2262}},
{{6'sd-27, 10'sd-261, 10'sd486}, {11'sd-803, 10'sd463, 8'sd-96}, {13'sd2816, 12'sd-1210, 12'sd1559}},
{{12'sd2011, 11'sd623, 10'sd346}, {12'sd-1605, 12'sd1158, 12'sd-1213}, {13'sd-3299, 12'sd1084, 13'sd-3038}},
{{9'sd-160, 10'sd258, 13'sd-2232}, {13'sd3413, 13'sd2610, 13'sd-2133}, {12'sd-1624, 11'sd538, 12'sd-1377}},
{{12'sd-1306, 12'sd1180, 10'sd-428}, {13'sd-2414, 11'sd695, 13'sd-2720}, {12'sd1793, 12'sd-1439, 11'sd630}},
{{9'sd-134, 7'sd40, 11'sd580}, {12'sd1959, 12'sd1639, 12'sd1189}, {11'sd536, 13'sd2937, 12'sd-1169}},
{{12'sd-1212, 13'sd-2949, 11'sd625}, {12'sd-1974, 13'sd2087, 11'sd-671}, {11'sd952, 11'sd-694, 11'sd526}},
{{12'sd1105, 7'sd61, 12'sd2007}, {13'sd-2165, 13'sd2399, 11'sd-948}, {8'sd70, 12'sd-1707, 13'sd2554}},
{{12'sd2020, 13'sd3118, 13'sd-2125}, {11'sd658, 11'sd625, 12'sd-1109}, {13'sd-2702, 10'sd-427, 12'sd1105}},
{{12'sd1362, 12'sd1745, 10'sd288}, {11'sd-848, 12'sd1835, 12'sd-1707}, {12'sd-1419, 12'sd1028, 12'sd-1601}},
{{12'sd-1405, 8'sd98, 10'sd326}, {13'sd-2541, 12'sd1733, 9'sd226}, {13'sd2279, 12'sd-1193, 10'sd434}},
{{13'sd3024, 12'sd1588, 12'sd1625}, {13'sd-3012, 8'sd93, 9'sd-214}, {13'sd-2167, 12'sd1325, 8'sd-77}},
{{12'sd1350, 9'sd-173, 12'sd1088}, {13'sd-3108, 12'sd-1716, 12'sd1874}, {13'sd2194, 10'sd-365, 12'sd1513}},
{{12'sd-1253, 13'sd2703, 12'sd1883}, {12'sd1080, 13'sd2586, 12'sd-1778}, {10'sd-438, 8'sd89, 8'sd93}},
{{12'sd1459, 8'sd127, 11'sd814}, {13'sd-2368, 12'sd-1865, 12'sd1587}, {9'sd-245, 12'sd-1549, 11'sd652}},
{{9'sd-253, 13'sd-2352, 13'sd2164}, {12'sd-1697, 10'sd261, 11'sd675}, {13'sd-2441, 12'sd1916, 12'sd-1039}},
{{11'sd585, 12'sd1767, 12'sd1594}, {10'sd-298, 11'sd-842, 13'sd2349}, {12'sd-1562, 12'sd1465, 13'sd3755}},
{{10'sd350, 11'sd-605, 11'sd828}, {10'sd345, 13'sd2204, 11'sd-829}, {13'sd2117, 10'sd-329, 12'sd1484}},
{{7'sd-33, 13'sd-2104, 9'sd-191}, {11'sd-721, 13'sd-3043, 10'sd-486}, {10'sd409, 12'sd-1709, 11'sd-940}},
{{13'sd2250, 13'sd-2293, 12'sd1318}, {12'sd1518, 9'sd-190, 13'sd-2143}, {12'sd-1237, 11'sd-668, 12'sd-1555}},
{{13'sd2244, 12'sd-1103, 11'sd-769}, {12'sd-1128, 12'sd1031, 13'sd-2526}, {13'sd-2656, 13'sd-2160, 12'sd-1867}},
{{12'sd1133, 11'sd862, 13'sd-2312}, {12'sd-1197, 12'sd1945, 11'sd-539}, {13'sd-2371, 12'sd-1792, 11'sd584}},
{{10'sd-491, 13'sd-2239, 13'sd2327}, {12'sd-1588, 12'sd1851, 12'sd2008}, {12'sd-1264, 13'sd2534, 12'sd1571}},
{{12'sd1620, 12'sd1843, 13'sd2574}, {9'sd-149, 12'sd1955, 11'sd905}, {13'sd-2099, 12'sd-1108, 12'sd1928}},
{{11'sd520, 13'sd2368, 12'sd1931}, {10'sd-287, 10'sd290, 12'sd1215}, {12'sd1085, 10'sd-279, 11'sd-790}},
{{13'sd-2494, 13'sd2130, 13'sd-2871}, {12'sd-1831, 11'sd-604, 12'sd1731}, {9'sd-223, 11'sd899, 13'sd-2220}},
{{9'sd-224, 13'sd-2253, 12'sd-1561}, {12'sd-1727, 12'sd1522, 12'sd-1578}, {11'sd-985, 12'sd1412, 10'sd426}},
{{12'sd-1999, 11'sd-927, 12'sd-1149}, {12'sd-1985, 12'sd1774, 8'sd87}, {12'sd-1600, 13'sd-2436, 11'sd-840}}},
{
{{9'sd190, 13'sd2351, 13'sd2825}, {13'sd2960, 13'sd2743, 11'sd-881}, {12'sd-1706, 11'sd-887, 11'sd-994}},
{{12'sd-2000, 10'sd-344, 13'sd-2056}, {12'sd-1668, 13'sd2816, 11'sd-603}, {11'sd873, 13'sd2644, 13'sd2256}},
{{10'sd385, 12'sd-1524, 12'sd1334}, {13'sd-2824, 13'sd2322, 12'sd1683}, {12'sd-1826, 13'sd-2923, 12'sd1628}},
{{12'sd-1032, 11'sd855, 12'sd-1914}, {12'sd2035, 11'sd923, 12'sd2002}, {13'sd-3128, 13'sd-2173, 11'sd548}},
{{11'sd777, 12'sd1930, 12'sd1473}, {11'sd1020, 11'sd-942, 11'sd513}, {13'sd2141, 12'sd1392, 7'sd43}},
{{12'sd1486, 11'sd926, 13'sd-2122}, {8'sd-112, 13'sd2670, 12'sd1384}, {11'sd-774, 13'sd-2306, 12'sd1454}},
{{9'sd238, 11'sd651, 13'sd2678}, {12'sd-1588, 11'sd-855, 9'sd174}, {11'sd-538, 11'sd824, 9'sd-161}},
{{10'sd364, 13'sd2133, 13'sd-3396}, {13'sd-2616, 10'sd294, 10'sd480}, {13'sd2796, 13'sd2628, 8'sd-103}},
{{8'sd98, 11'sd564, 12'sd1088}, {12'sd-1588, 11'sd584, 12'sd1853}, {11'sd851, 10'sd509, 13'sd-2230}},
{{11'sd521, 13'sd2982, 11'sd-745}, {12'sd1486, 12'sd1190, 13'sd-2552}, {13'sd-2841, 12'sd-1128, 11'sd545}},
{{13'sd-3585, 13'sd-3602, 12'sd1789}, {9'sd-184, 12'sd1920, 13'sd-2954}, {12'sd-1282, 13'sd-2240, 11'sd907}},
{{11'sd-996, 13'sd-2564, 9'sd-179}, {11'sd789, 12'sd-1050, 13'sd-2712}, {9'sd181, 12'sd-1662, 10'sd445}},
{{12'sd1692, 9'sd-163, 12'sd-1214}, {12'sd-1741, 13'sd-2343, 13'sd-2441}, {6'sd30, 13'sd-2277, 13'sd-2772}},
{{11'sd610, 13'sd-2795, 13'sd2967}, {13'sd-2634, 4'sd4, 8'sd115}, {10'sd321, 12'sd-1719, 12'sd1614}},
{{14'sd4173, 12'sd1729, 13'sd-2686}, {12'sd-1061, 11'sd-1016, 13'sd-3537}, {10'sd-457, 13'sd2590, 12'sd-1034}},
{{12'sd1806, 12'sd1576, 13'sd-3390}, {12'sd-1154, 13'sd2086, 11'sd732}, {12'sd1048, 12'sd1504, 12'sd-1301}},
{{13'sd-2845, 10'sd380, 10'sd-452}, {13'sd2225, 11'sd587, 12'sd-1431}, {10'sd-303, 12'sd1863, 12'sd1894}},
{{13'sd3459, 13'sd2486, 11'sd-857}, {10'sd-395, 10'sd264, 13'sd2065}, {13'sd2906, 11'sd-818, 8'sd-106}},
{{13'sd3045, 11'sd-1018, 13'sd2224}, {12'sd-1192, 12'sd-1104, 13'sd2745}, {12'sd1519, 12'sd1750, 11'sd641}},
{{13'sd-2089, 5'sd-12, 11'sd757}, {13'sd-2495, 12'sd1203, 11'sd-1002}, {12'sd1704, 11'sd905, 10'sd-299}},
{{12'sd2023, 12'sd1566, 11'sd-775}, {13'sd-2067, 10'sd503, 13'sd-2484}, {12'sd1313, 13'sd2521, 13'sd-2387}},
{{12'sd1622, 10'sd-504, 12'sd-1784}, {11'sd-716, 13'sd-3345, 11'sd-657}, {13'sd2741, 13'sd2068, 12'sd2035}},
{{12'sd-1040, 12'sd1662, 13'sd-2693}, {12'sd-2004, 13'sd-2986, 13'sd-3065}, {12'sd-1426, 11'sd683, 11'sd878}},
{{9'sd-141, 12'sd1981, 12'sd1297}, {13'sd-2262, 13'sd-2869, 12'sd-1384}, {11'sd878, 12'sd-1764, 10'sd-373}},
{{12'sd-1221, 12'sd-1882, 12'sd-1314}, {12'sd-1142, 13'sd2807, 13'sd2159}, {13'sd-2316, 10'sd-297, 11'sd553}},
{{9'sd219, 13'sd2485, 10'sd-424}, {12'sd1670, 13'sd2258, 13'sd-2552}, {13'sd-3539, 13'sd2255, 13'sd-3165}},
{{10'sd375, 12'sd-1387, 8'sd-92}, {13'sd-2896, 12'sd1964, 13'sd-2712}, {13'sd-2626, 11'sd-999, 13'sd-2844}},
{{12'sd1493, 13'sd-2302, 13'sd-2050}, {8'sd-89, 11'sd-852, 13'sd2182}, {12'sd-1744, 11'sd-650, 13'sd3673}},
{{13'sd-2169, 13'sd2215, 13'sd2118}, {11'sd585, 13'sd-2592, 12'sd-1645}, {11'sd-625, 11'sd888, 12'sd-1262}},
{{12'sd1526, 12'sd1903, 12'sd1933}, {7'sd-41, 13'sd-2290, 12'sd1138}, {12'sd1089, 8'sd76, 13'sd-2480}},
{{12'sd1596, 13'sd-2809, 13'sd-2158}, {13'sd2945, 12'sd1941, 11'sd608}, {13'sd-2057, 8'sd-92, 13'sd-2524}},
{{12'sd1389, 13'sd-2188, 13'sd-2372}, {9'sd211, 12'sd-1152, 11'sd692}, {13'sd3493, 12'sd1215, 11'sd-664}},
{{10'sd269, 11'sd-705, 12'sd1418}, {12'sd-1674, 11'sd-951, 13'sd-2825}, {11'sd632, 11'sd-554, 8'sd64}},
{{12'sd1121, 12'sd1220, 13'sd3154}, {12'sd-1369, 13'sd2097, 11'sd842}, {12'sd1188, 12'sd-1624, 12'sd1166}},
{{12'sd1870, 13'sd2779, 13'sd-2995}, {11'sd934, 12'sd-1191, 11'sd945}, {10'sd-376, 13'sd-2224, 11'sd-753}},
{{12'sd-1710, 11'sd597, 9'sd-232}, {12'sd1748, 12'sd-1983, 13'sd3069}, {12'sd1794, 13'sd2143, 12'sd-1250}},
{{13'sd-2063, 12'sd-1203, 12'sd1230}, {13'sd2646, 12'sd-1238, 8'sd-95}, {11'sd-706, 11'sd609, 13'sd3162}},
{{11'sd769, 11'sd-873, 11'sd-693}, {13'sd2268, 13'sd2749, 11'sd927}, {13'sd2632, 11'sd761, 12'sd-1734}},
{{13'sd2213, 12'sd-1764, 13'sd2076}, {9'sd155, 12'sd1746, 13'sd-2167}, {13'sd-2622, 7'sd40, 10'sd307}},
{{9'sd-185, 13'sd-2965, 12'sd-1757}, {12'sd1612, 7'sd-52, 10'sd478}, {11'sd567, 12'sd1232, 12'sd-1512}},
{{13'sd2808, 13'sd2315, 12'sd-1512}, {13'sd-2472, 9'sd223, 13'sd-2969}, {10'sd331, 12'sd1460, 11'sd716}},
{{12'sd1632, 13'sd2982, 11'sd857}, {10'sd470, 11'sd-977, 12'sd1897}, {12'sd-1429, 11'sd-865, 12'sd-1930}},
{{12'sd-1675, 12'sd-1568, 13'sd-2232}, {11'sd-769, 12'sd-1199, 8'sd-69}, {11'sd-662, 8'sd125, 13'sd-2851}},
{{11'sd615, 10'sd-363, 11'sd813}, {12'sd-1208, 11'sd-738, 12'sd-1466}, {12'sd-1099, 11'sd-1001, 12'sd1218}},
{{13'sd2963, 13'sd-2377, 12'sd1873}, {12'sd-1377, 12'sd1083, 12'sd-1551}, {13'sd-2377, 11'sd-718, 11'sd715}},
{{10'sd495, 11'sd814, 12'sd-1442}, {12'sd1196, 11'sd536, 10'sd505}, {13'sd-2237, 12'sd-1031, 11'sd617}},
{{11'sd-903, 13'sd2488, 13'sd2456}, {12'sd1360, 12'sd1762, 12'sd-1930}, {13'sd2181, 9'sd-130, 12'sd-1115}},
{{11'sd963, 12'sd-1579, 7'sd-41}, {12'sd1742, 12'sd1151, 13'sd-3022}, {11'sd-659, 12'sd1726, 12'sd-1360}},
{{13'sd-2478, 12'sd-1603, 11'sd-602}, {12'sd-1064, 13'sd2684, 11'sd-861}, {11'sd-679, 10'sd266, 11'sd-678}},
{{12'sd-1141, 12'sd1174, 11'sd-559}, {13'sd-2303, 12'sd2034, 13'sd2075}, {12'sd1180, 12'sd1727, 10'sd420}},
{{10'sd276, 12'sd1819, 13'sd-2372}, {12'sd1108, 12'sd1282, 12'sd1800}, {10'sd410, 10'sd-485, 13'sd-3204}},
{{8'sd-67, 12'sd1078, 12'sd-1143}, {12'sd-1965, 13'sd2328, 12'sd2046}, {12'sd-2033, 12'sd1981, 13'sd-2844}},
{{13'sd-2463, 12'sd1432, 13'sd2806}, {13'sd-2117, 13'sd2183, 10'sd-347}, {14'sd-4141, 13'sd2189, 12'sd-2045}},
{{11'sd-647, 12'sd1650, 11'sd-601}, {12'sd-1603, 12'sd1117, 13'sd-2453}, {11'sd730, 13'sd2122, 8'sd100}},
{{11'sd-977, 12'sd1334, 12'sd-1719}, {13'sd-2927, 13'sd-2961, 10'sd-306}, {12'sd-1114, 11'sd703, 10'sd362}},
{{12'sd1111, 13'sd-2563, 11'sd-808}, {11'sd-992, 12'sd1067, 13'sd2058}, {12'sd-1578, 12'sd-2030, 12'sd1249}},
{{11'sd-951, 13'sd-2753, 13'sd-2819}, {11'sd-554, 11'sd-551, 12'sd1129}, {9'sd217, 12'sd1334, 7'sd61}},
{{10'sd-361, 12'sd-1399, 13'sd-2254}, {12'sd-2040, 12'sd-2018, 11'sd747}, {9'sd-215, 12'sd-1678, 10'sd-386}},
{{10'sd-381, 10'sd-359, 11'sd588}, {9'sd-180, 12'sd-1115, 11'sd-688}, {11'sd-758, 11'sd-560, 13'sd2215}},
{{13'sd2467, 12'sd1843, 10'sd495}, {11'sd987, 9'sd-223, 13'sd2069}, {13'sd-2095, 13'sd-2563, 12'sd2016}},
{{12'sd-1142, 10'sd-511, 12'sd-1850}, {13'sd2688, 12'sd1036, 12'sd-1444}, {13'sd-2503, 11'sd-951, 12'sd1303}},
{{11'sd-725, 13'sd-2356, 11'sd-940}, {13'sd-2200, 12'sd1976, 11'sd-582}, {13'sd-2168, 12'sd-1584, 8'sd-117}},
{{10'sd317, 10'sd-472, 13'sd-2275}, {13'sd-2963, 13'sd-2067, 10'sd-334}, {11'sd-852, 11'sd1019, 12'sd1111}},
{{12'sd-2023, 9'sd186, 10'sd418}, {11'sd-787, 8'sd-98, 11'sd-1002}, {13'sd-2609, 12'sd-1854, 10'sd375}}},
{
{{12'sd1045, 11'sd676, 13'sd2649}, {13'sd2380, 11'sd827, 10'sd-378}, {10'sd-291, 12'sd1924, 12'sd-1211}},
{{12'sd1517, 12'sd-1304, 12'sd-1340}, {12'sd1838, 11'sd-667, 8'sd-121}, {13'sd2689, 12'sd-1149, 7'sd58}},
{{12'sd-1103, 10'sd-311, 13'sd-2545}, {12'sd-1770, 8'sd108, 13'sd2619}, {11'sd729, 12'sd1486, 12'sd1342}},
{{12'sd1418, 13'sd-2731, 13'sd-3043}, {13'sd2631, 10'sd489, 9'sd-231}, {12'sd1612, 11'sd-1005, 12'sd1281}},
{{13'sd3136, 12'sd1096, 10'sd-371}, {7'sd41, 9'sd238, 12'sd-1601}, {11'sd789, 12'sd-1800, 13'sd2599}},
{{11'sd820, 13'sd-2878, 13'sd-2153}, {11'sd984, 9'sd-172, 10'sd-423}, {11'sd-769, 11'sd-595, 11'sd1013}},
{{11'sd577, 10'sd413, 11'sd-744}, {11'sd-988, 12'sd-1251, 13'sd2409}, {12'sd-1081, 13'sd2711, 12'sd-1622}},
{{13'sd2150, 11'sd-699, 10'sd-345}, {13'sd2242, 8'sd127, 13'sd-2544}, {10'sd472, 12'sd-1793, 13'sd2284}},
{{12'sd-1071, 12'sd1707, 12'sd1495}, {12'sd1779, 11'sd-642, 8'sd-111}, {10'sd-313, 12'sd1061, 10'sd-257}},
{{12'sd2047, 12'sd1381, 12'sd-1793}, {12'sd1370, 12'sd-1976, 12'sd1345}, {12'sd-1083, 8'sd-120, 13'sd2657}},
{{13'sd-3364, 11'sd-751, 13'sd-2662}, {10'sd262, 9'sd-200, 12'sd1778}, {12'sd-1091, 12'sd1960, 11'sd739}},
{{11'sd981, 12'sd-1686, 12'sd1997}, {13'sd-2699, 12'sd1427, 13'sd-2969}, {8'sd-93, 12'sd-1803, 11'sd609}},
{{13'sd-2977, 13'sd-2539, 13'sd-2317}, {13'sd-2759, 13'sd-2221, 12'sd-1079}, {10'sd-353, 13'sd-2634, 13'sd2529}},
{{12'sd-1812, 8'sd110, 11'sd-621}, {10'sd-414, 12'sd1368, 13'sd2203}, {12'sd-1360, 13'sd-2070, 13'sd2423}},
{{13'sd2700, 11'sd-881, 13'sd-3384}, {12'sd-1352, 12'sd2037, 13'sd-2111}, {13'sd2593, 10'sd-274, 10'sd-361}},
{{13'sd2331, 8'sd64, 13'sd-2760}, {11'sd913, 12'sd1102, 10'sd-485}, {12'sd1974, 13'sd2890, 11'sd-606}},
{{12'sd1240, 11'sd842, 12'sd-1039}, {12'sd1604, 13'sd-2550, 12'sd-1188}, {13'sd2239, 13'sd2161, 12'sd1550}},
{{10'sd486, 10'sd293, 12'sd-1188}, {9'sd200, 12'sd1473, 12'sd-1295}, {13'sd2491, 13'sd2727, 11'sd912}},
{{10'sd283, 11'sd549, 12'sd-1661}, {12'sd-1385, 13'sd-2501, 12'sd-1192}, {13'sd2157, 12'sd1366, 13'sd2650}},
{{12'sd1158, 12'sd-1907, 11'sd-845}, {11'sd-598, 13'sd3154, 13'sd-2125}, {11'sd590, 12'sd-1747, 12'sd1442}},
{{13'sd2197, 12'sd1690, 12'sd-1376}, {13'sd-3339, 11'sd-940, 10'sd329}, {13'sd-2289, 13'sd2428, 10'sd287}},
{{12'sd1347, 12'sd1791, 13'sd-3592}, {11'sd524, 12'sd1713, 12'sd-1754}, {12'sd-1621, 12'sd1689, 11'sd-805}},
{{10'sd462, 13'sd-3524, 11'sd937}, {12'sd-1300, 13'sd-2730, 13'sd-2125}, {12'sd-1247, 12'sd-1628, 11'sd663}},
{{12'sd-2016, 12'sd-1816, 13'sd-3647}, {13'sd-2754, 12'sd1800, 9'sd141}, {9'sd151, 11'sd-581, 12'sd-1572}},
{{12'sd1905, 11'sd787, 13'sd3643}, {13'sd2383, 12'sd-1389, 12'sd-1871}, {13'sd-2331, 8'sd-84, 11'sd-954}},
{{12'sd1497, 12'sd-1453, 11'sd996}, {11'sd665, 11'sd1013, 13'sd-2808}, {11'sd948, 12'sd1244, 12'sd1224}},
{{13'sd-2512, 11'sd-518, 13'sd-2527}, {13'sd2326, 9'sd-204, 12'sd-1457}, {10'sd-489, 10'sd-275, 12'sd-1804}},
{{13'sd2316, 11'sd-849, 11'sd757}, {11'sd-595, 9'sd179, 11'sd791}, {10'sd272, 13'sd-3169, 13'sd-2507}},
{{12'sd-1668, 12'sd-1552, 13'sd-2048}, {12'sd1043, 9'sd143, 13'sd-2454}, {8'sd-116, 12'sd-1578, 13'sd2295}},
{{12'sd-1389, 8'sd-91, 8'sd67}, {7'sd33, 12'sd1548, 11'sd-581}, {9'sd-232, 13'sd3002, 12'sd1681}},
{{12'sd-2014, 9'sd195, 13'sd3129}, {10'sd498, 11'sd689, 12'sd-1177}, {13'sd2155, 11'sd-789, 9'sd-201}},
{{11'sd746, 13'sd-2189, 13'sd2949}, {12'sd-1609, 12'sd-1629, 11'sd618}, {11'sd831, 12'sd1562, 12'sd1209}},
{{12'sd-1632, 13'sd-2824, 10'sd-296}, {13'sd-2088, 11'sd-735, 13'sd-2569}, {13'sd-2254, 11'sd866, 10'sd-511}},
{{12'sd-1190, 12'sd-1887, 13'sd-2473}, {12'sd1380, 13'sd2055, 12'sd1779}, {11'sd-862, 12'sd-1404, 13'sd2483}},
{{13'sd3798, 10'sd507, 11'sd860}, {13'sd4077, 10'sd-440, 9'sd174}, {7'sd-61, 14'sd-5142, 14'sd-6269}},
{{13'sd-2183, 13'sd-2383, 12'sd-1722}, {13'sd2302, 13'sd-2936, 12'sd1708}, {10'sd-502, 13'sd-3145, 13'sd3171}},
{{12'sd1735, 12'sd1519, 13'sd2953}, {13'sd-2159, 12'sd1203, 12'sd-1910}, {9'sd-249, 13'sd2224, 12'sd1884}},
{{13'sd-2178, 13'sd2588, 12'sd-1571}, {11'sd-817, 12'sd1975, 13'sd2544}, {11'sd567, 11'sd1000, 12'sd-1060}},
{{7'sd-41, 10'sd-341, 12'sd-1148}, {12'sd-1751, 12'sd1444, 13'sd-2125}, {12'sd1661, 13'sd2562, 12'sd1341}},
{{12'sd1365, 8'sd-98, 11'sd891}, {12'sd-2020, 10'sd270, 13'sd3412}, {13'sd-3603, 9'sd204, 11'sd-774}},
{{12'sd2002, 12'sd-1349, 13'sd-2804}, {10'sd436, 12'sd1146, 9'sd-233}, {13'sd2864, 7'sd-37, 9'sd173}},
{{13'sd2622, 11'sd-778, 9'sd249}, {11'sd-580, 11'sd649, 13'sd-2051}, {10'sd486, 13'sd2537, 11'sd-628}},
{{13'sd-2873, 12'sd-1387, 11'sd845}, {7'sd32, 13'sd2624, 12'sd1335}, {12'sd1574, 10'sd387, 13'sd3297}},
{{11'sd-925, 10'sd-371, 12'sd-1979}, {12'sd-1481, 12'sd1792, 12'sd1722}, {8'sd-117, 11'sd755, 11'sd-608}},
{{11'sd-875, 12'sd1366, 12'sd1046}, {12'sd1775, 10'sd472, 12'sd1590}, {13'sd-2665, 13'sd-3155, 12'sd1177}},
{{11'sd923, 13'sd-3122, 13'sd2169}, {10'sd327, 10'sd485, 13'sd2276}, {13'sd-3159, 11'sd653, 13'sd-2369}},
{{13'sd2891, 12'sd-1147, 13'sd-2146}, {7'sd-36, 12'sd1857, 13'sd2100}, {9'sd-182, 12'sd1548, 9'sd-186}},
{{12'sd-1306, 12'sd-1239, 13'sd2983}, {11'sd-544, 11'sd-943, 11'sd-683}, {13'sd2487, 11'sd-549, 12'sd-1471}},
{{12'sd-1399, 12'sd-1830, 12'sd-1963}, {10'sd-260, 12'sd1838, 13'sd2189}, {12'sd1097, 12'sd-1983, 11'sd837}},
{{11'sd-832, 7'sd52, 13'sd2507}, {12'sd-1307, 12'sd1701, 13'sd2365}, {12'sd-1034, 13'sd-2903, 11'sd-704}},
{{12'sd-1287, 12'sd-1535, 12'sd-1331}, {13'sd-2279, 12'sd-1613, 13'sd2377}, {11'sd742, 10'sd-272, 13'sd3400}},
{{13'sd2469, 11'sd572, 10'sd-469}, {12'sd-1636, 8'sd-88, 12'sd-1922}, {12'sd1563, 10'sd392, 11'sd729}},
{{13'sd-3738, 10'sd-352, 13'sd2259}, {12'sd1411, 12'sd-1084, 8'sd-81}, {13'sd-2747, 12'sd-1466, 10'sd-366}},
{{13'sd-2335, 11'sd-937, 13'sd-2135}, {13'sd-2945, 11'sd547, 12'sd1907}, {13'sd2410, 12'sd1538, 12'sd1346}},
{{12'sd-1271, 9'sd-182, 12'sd1910}, {11'sd-717, 10'sd327, 11'sd974}, {13'sd2203, 12'sd2039, 11'sd-998}},
{{12'sd1209, 13'sd-2363, 9'sd-163}, {13'sd-2831, 12'sd-1312, 11'sd-975}, {13'sd-3065, 13'sd-2852, 11'sd-849}},
{{11'sd-576, 8'sd87, 13'sd-2142}, {11'sd828, 10'sd-445, 12'sd-1674}, {12'sd-1665, 10'sd336, 11'sd-656}},
{{12'sd1224, 12'sd1441, 8'sd121}, {12'sd1863, 12'sd1902, 12'sd-1446}, {13'sd2331, 10'sd329, 12'sd-1423}},
{{11'sd546, 12'sd1604, 9'sd-170}, {11'sd-901, 12'sd-1386, 13'sd-2614}, {11'sd858, 12'sd-1652, 10'sd397}},
{{12'sd1592, 13'sd2244, 11'sd581}, {13'sd2457, 12'sd-1131, 10'sd-259}, {12'sd1430, 12'sd-1740, 12'sd1097}},
{{13'sd2368, 12'sd1966, 12'sd1026}, {11'sd-524, 12'sd1553, 11'sd981}, {11'sd1019, 12'sd-1457, 13'sd2428}},
{{10'sd-405, 13'sd-3052, 12'sd-1398}, {13'sd-2929, 11'sd829, 12'sd-1054}, {13'sd-2120, 13'sd2432, 12'sd1071}},
{{12'sd1880, 12'sd-1865, 12'sd1156}, {11'sd-937, 9'sd-232, 13'sd-2447}, {13'sd-2093, 12'sd-1182, 11'sd-838}},
{{11'sd764, 11'sd-863, 12'sd-1709}, {10'sd-371, 13'sd-2474, 13'sd-2883}, {13'sd2314, 12'sd-1353, 13'sd-2599}}}}};


// 2D Register to store convolution biases: [ConvLayer][Bias]
// Fixed-point format: 16 fractional bits
reg signed [31:0] conv_biases[0:4][0:63] = '{
// Biases for conv1_bias
{
  14'sd7150,
  14'sd7533,
  15'sd11206,
  15'sd-11033,
  14'sd-6885,
  12'sd2030,
  13'sd-3330,
  15'sd-8258,
  14'sd7971,
  15'sd-9152,
  12'sd1472,
  15'sd10162,
  13'sd-2538,
  15'sd-9351,
  14'sd-4750,
  13'sd3784,
  14'sd-7951,
  15'sd-11688,
  15'sd-11214,
  14'sd-4997,
  14'sd-5132,
  15'sd-10462,
  15'sd-9103,
  14'sd-5330,
  15'sd-10393,
  14'sd6746,
  1'sd0,
  13'sd2248,
  13'sd-3264,
  14'sd7197,
  15'sd-9150,
  14'sd5167,
  14'sd-7213,
  14'sd6323,
  12'sd1093,
  14'sd-4811,
  14'sd7308,
  15'sd-8254,
  14'sd-6724,
  15'sd9698,
  15'sd-8239,
  12'sd-1831,
  14'sd-4773,
  12'sd-1583,
  15'sd10951,
  14'sd-4633,
  14'sd6288,
  14'sd-6338,
  15'sd9657,
  13'sd3758,
  14'sd-5005,
  15'sd9179,
  9'sd-213,
  14'sd-6278,
  14'sd-6562,
  10'sd307,
  14'sd-4219,
  12'sd-1221,
  15'sd10295,
  12'sd-1400,
  15'sd-11286,
  12'sd1961,
  10'sd382,
  4'sd-6
},
// Biases for conv2_bias
{
  10'sd493,
  13'sd-2052,
  13'sd2083,
  12'sd1764,
  12'sd-1862,
  11'sd-669,
  12'sd1089,
  12'sd1489,
  13'sd-2172,
  12'sd1353,
  12'sd-1545,
  12'sd1739,
  13'sd-2834,
  12'sd2046,
  12'sd-1094,
  12'sd1356,
  9'sd-184,
  10'sd324,
  12'sd-1397,
  13'sd-2491,
  12'sd1239,
  9'sd218,
  12'sd-1833,
  13'sd2357,
  10'sd-357,
  9'sd201,
  11'sd-560,
  7'sd55,
  11'sd-996,
  11'sd808,
  10'sd-462,
  12'sd-1352,
  12'sd1349,
  10'sd281,
  13'sd2290,
  12'sd1240,
  12'sd1578,
  13'sd2224,
  10'sd-474,
  13'sd2061,
  13'sd-2242,
  12'sd1972,
  12'sd1826,
  10'sd-420,
  8'sd-90,
  12'sd1405,
  8'sd109,
  12'sd1239,
  9'sd180,
  11'sd810,
  5'sd9,
  12'sd1981,
  12'sd-1545,
  4'sd-7,
  12'sd-1689,
  11'sd995,
  11'sd602,
  12'sd-1316,
  13'sd2961,
  13'sd2694,
  10'sd-473,
  11'sd852,
  10'sd-257,
  11'sd-855
},
// Biases for conv3_bias
{
  12'sd-1383,
  12'sd-1827,
  12'sd1734,
  12'sd1519,
  13'sd-2296,
  10'sd319,
  13'sd-2551,
  13'sd-2773,
  12'sd2025,
  12'sd1065,
  13'sd3145,
  12'sd1237,
  13'sd2219,
  12'sd1538,
  13'sd2084,
  13'sd2694,
  5'sd-10,
  12'sd1086,
  10'sd-357,
  13'sd3017,
  12'sd-1837,
  9'sd-210,
  11'sd780,
  13'sd-3065,
  13'sd2617,
  13'sd2897,
  13'sd-3364,
  12'sd1877,
  12'sd1372,
  13'sd3160,
  12'sd1704,
  13'sd-3477,
  13'sd-2783,
  13'sd2811,
  13'sd-2195,
  13'sd2893,
  13'sd-2185,
  13'sd2500,
  8'sd-70,
  8'sd104,
  12'sd-1247,
  12'sd-2001,
  12'sd2047,
  12'sd1359,
  13'sd-3002,
  13'sd2389,
  12'sd1339,
  10'sd447,
  11'sd-951,
  11'sd-703,
  12'sd-1688,
  11'sd558,
  13'sd-2063,
  13'sd-2126,
  11'sd-664,
  12'sd1255,
  13'sd2456,
  12'sd1258,
  12'sd1683,
  12'sd1286,
  13'sd-3082,
  12'sd1111,
  12'sd1820,
  10'sd-334
},
// Biases for conv4_bias
{
  14'sd4183,
  14'sd4191,
  7'sd45,
  12'sd1035,
  13'sd3535,
  10'sd-463,
  13'sd2307,
  13'sd4094,
  9'sd149,
  11'sd529,
  13'sd-3700,
  13'sd-2589,
  8'sd-111,
  13'sd-2766,
  11'sd672,
  10'sd-490,
  11'sd636,
  13'sd2981,
  13'sd3413,
  8'sd83,
  10'sd321,
  11'sd-904,
  12'sd-1905,
  13'sd-2767,
  9'sd-244,
  12'sd1413,
  13'sd-3590,
  13'sd-2389,
  12'sd-1828,
  13'sd3174,
  12'sd1900,
  10'sd358,
  12'sd-1384,
  14'sd4129,
  12'sd-1757,
  13'sd3050,
  13'sd2615,
  13'sd4004,
  11'sd-949,
  12'sd-1030,
  10'sd-290,
  13'sd2824,
  13'sd-2182,
  12'sd1123,
  8'sd123,
  10'sd-258,
  8'sd66,
  10'sd424,
  10'sd510,
  9'sd240,
  13'sd-2070,
  10'sd417,
  11'sd-965,
  11'sd535,
  13'sd-2618,
  10'sd-370,
  13'sd-2924,
  12'sd-1630,
  9'sd-193,
  11'sd-991,
  12'sd1309,
  10'sd342,
  14'sd-4137,
  13'sd-2225
},
// Biases for conv5_bias
{
  12'sd1388,
  13'sd2049,
  12'sd1099
}};
initial begin
    Weights = conv_weights
    Biases = conv_biases
end


endmodule